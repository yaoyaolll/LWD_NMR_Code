library verilog;
use verilog.vl_types.all;
entity off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_3 is
    port(
        i_6             : in     vl_logic_vector(1 downto 1);
        i_7             : in     vl_logic_vector(0 downto 0);
        GLA             : in     vl_logic;
        DUMP_0_dump_on  : out    vl_logic;
        off_on_state_1_state_over: out    vl_logic;
        state1ms_choice_0_reset_out: in     vl_logic
    );
end off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_3;
