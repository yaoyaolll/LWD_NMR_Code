`timescale 1 ns/100 ps
// Version: v11.9 SP6 11.9.6.7
// File used only for Simulation


module PLLBA(
       CLKA,
       EXTFB,
       POWERDOWN,
       GLA,
       LOCK,
       GLB,
       YB,
       GLC,
       YC,
       OADIV0,
       OADIV1,
       OADIV2,
       OADIV3,
       OADIV4,
       OAMUX0,
       OAMUX1,
       OAMUX2,
       DLYGLA0,
       DLYGLA1,
       DLYGLA2,
       DLYGLA3,
       DLYGLA4,
       OBDIV0,
       OBDIV1,
       OBDIV2,
       OBDIV3,
       OBDIV4,
       OBMUX0,
       OBMUX1,
       OBMUX2,
       DLYYB0,
       DLYYB1,
       DLYYB2,
       DLYYB3,
       DLYYB4,
       DLYGLB0,
       DLYGLB1,
       DLYGLB2,
       DLYGLB3,
       DLYGLB4,
       OCDIV0,
       OCDIV1,
       OCDIV2,
       OCDIV3,
       OCDIV4,
       OCMUX0,
       OCMUX1,
       OCMUX2,
       DLYYC0,
       DLYYC1,
       DLYYC2,
       DLYYC3,
       DLYYC4,
       DLYGLC0,
       DLYGLC1,
       DLYGLC2,
       DLYGLC3,
       DLYGLC4,
       FINDIV0,
       FINDIV1,
       FINDIV2,
       FINDIV3,
       FINDIV4,
       FINDIV5,
       FINDIV6,
       FBDIV0,
       FBDIV1,
       FBDIV2,
       FBDIV3,
       FBDIV4,
       FBDIV5,
       FBDIV6,
       FBDLY0,
       FBDLY1,
       FBDLY2,
       FBDLY3,
       FBDLY4,
       FBSEL0,
       FBSEL1,
       XDLYSEL,
       VCOSEL0,
       VCOSEL1,
       VCOSEL2
    );
input  CLKA;
input  EXTFB;
input  POWERDOWN;
output GLA;
output LOCK;
output GLB;
output YB;
output GLC;
output YC;
input  OADIV0;
input  OADIV1;
input  OADIV2;
input  OADIV3;
input  OADIV4;
input  OAMUX0;
input  OAMUX1;
input  OAMUX2;
input  DLYGLA0;
input  DLYGLA1;
input  DLYGLA2;
input  DLYGLA3;
input  DLYGLA4;
input  OBDIV0;
input  OBDIV1;
input  OBDIV2;
input  OBDIV3;
input  OBDIV4;
input  OBMUX0;
input  OBMUX1;
input  OBMUX2;
input  DLYYB0;
input  DLYYB1;
input  DLYYB2;
input  DLYYB3;
input  DLYYB4;
input  DLYGLB0;
input  DLYGLB1;
input  DLYGLB2;
input  DLYGLB3;
input  DLYGLB4;
input  OCDIV0;
input  OCDIV1;
input  OCDIV2;
input  OCDIV3;
input  OCDIV4;
input  OCMUX0;
input  OCMUX1;
input  OCMUX2;
input  DLYYC0;
input  DLYYC1;
input  DLYYC2;
input  DLYYC3;
input  DLYYC4;
input  DLYGLC0;
input  DLYGLC1;
input  DLYGLC2;
input  DLYGLC3;
input  DLYGLC4;
input  FINDIV0;
input  FINDIV1;
input  FINDIV2;
input  FINDIV3;
input  FINDIV4;
input  FINDIV5;
input  FINDIV6;
input  FBDIV0;
input  FBDIV1;
input  FBDIV2;
input  FBDIV3;
input  FBDIV4;
input  FBDIV5;
input  FBDIV6;
input  FBDLY0;
input  FBDLY1;
input  FBDLY2;
input  FBDLY3;
input  FBDLY4;
input  FBSEL0;
input  FBSEL1;
input  XDLYSEL;
input  VCOSEL0;
input  VCOSEL1;
input  VCOSEL2;

    wire GND, SDOUT, FB, EXTFBDLY, GLADLY, LOCKDLY, GLBDLY, YBDLY, 
        GLCDLY, YCDLY, VCODLY;
    wire GND_power_net1;
    assign GND = GND_power_net1;
    
    PLL_SDF #( .VCOFREQUENCY(100.000000) )  pll_sdf_0 (.CLKA(CLKA), 
        .EXTFB(EXTFBDLY), .POWERDOWN(POWERDOWN), .GLAOUT(GLADLY), 
        .LOCKOUT(LOCKDLY), .GLBOUT(GLBDLY), .YBOUT(YBDLY), .GLCOUT(
        GLCDLY), .YCOUT(YCDLY), .OADIV0(OADIV0), .OADIV1(OADIV1), 
        .OADIV2(OADIV2), .OADIV3(OADIV3), .OADIV4(OADIV4), .OAMUX0(
        OAMUX0), .OAMUX1(OAMUX1), .OAMUX2(OAMUX2), .DLYGLA0(DLYGLA0), 
        .DLYGLA1(DLYGLA1), .DLYGLA2(DLYGLA2), .DLYGLA3(DLYGLA3), 
        .DLYGLA4(DLYGLA4), .OBDIV0(OBDIV0), .OBDIV1(OBDIV1), .OBDIV2(
        OBDIV2), .OBDIV3(OBDIV3), .OBDIV4(OBDIV4), .OBMUX0(OBMUX0), 
        .OBMUX1(OBMUX1), .OBMUX2(OBMUX2), .DLYYB0(DLYYB0), .DLYYB1(
        DLYYB1), .DLYYB2(DLYYB2), .DLYYB3(DLYYB3), .DLYYB4(DLYYB4), 
        .DLYGLB0(DLYGLB0), .DLYGLB1(DLYGLB1), .DLYGLB2(DLYGLB2), 
        .DLYGLB3(DLYGLB3), .DLYGLB4(DLYGLB4), .OCDIV0(OCDIV0), .OCDIV1(
        OCDIV1), .OCDIV2(OCDIV2), .OCDIV3(OCDIV3), .OCDIV4(OCDIV4), 
        .OCMUX0(OCMUX0), .OCMUX1(OCMUX1), .OCMUX2(OCMUX2), .DLYYC0(
        DLYYC0), .DLYYC1(DLYYC1), .DLYYC2(DLYYC2), .DLYYC3(DLYYC3), 
        .DLYYC4(DLYYC4), .DLYGLC0(DLYGLC0), .DLYGLC1(DLYGLC1), 
        .DLYGLC2(DLYGLC2), .DLYGLC3(DLYGLC3), .DLYGLC4(DLYGLC4), 
        .FINDIV0(FINDIV0), .FINDIV1(FINDIV1), .FINDIV2(FINDIV2), 
        .FINDIV3(FINDIV3), .FINDIV4(FINDIV4), .FINDIV5(FINDIV5), 
        .FINDIV6(FINDIV6), .FBDIV0(FBDIV0), .FBDIV1(FBDIV1), .FBDIV2(
        FBDIV2), .FBDIV3(FBDIV3), .FBDIV4(FBDIV4), .FBDIV5(FBDIV5), 
        .FBDIV6(FBDIV6), .FBDLY0(FBDLY0), .FBDLY1(FBDLY1), .FBDLY2(
        FBDLY2), .FBDLY3(FBDLY3), .FBDLY4(FBDLY4), .FBSEL0(FBSEL0), 
        .FBSEL1(FBSEL1), .XDLYSEL(XDLYSEL), .VCOSEL0(VCOSEL0), 
        .VCOSEL1(VCOSEL1), .VCOSEL2(VCOSEL2), .INTFB(FB), .VCOOUT(
        VCODLY));
    PLL_DLY_SDF #( .VCOFREQUENCY(100.000000) )  pll_dly_sdf_0 (.GLA(
        GLA), .LOCK(LOCK), .GLB(GLB), .YB(YB), .GLC(GLC), .YC(YC), 
        .GLAIN(GLADLY), .LOCKIN(LOCKDLY), .GLBIN(GLBDLY), .YBIN(YBDLY), 
        .GLCIN(GLCDLY), .YCIN(YCDLY), .EXTFBOUT(EXTFBDLY), .EXTFBIN(
        EXTFB), .VCOIN(VCODLY), .PLLOUT(FB));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module NMR_TOP(
       ADC,
       OCX40MHz,
       XRD,
       ddsclkout,
       gpio,
       tri_ctrl,
       xa,
       xwe,
       zcs2,
       Acq_clk,
       GLA,
       Q1Q8,
       Q2Q7,
       Q3Q6,
       Q4Q5,
       cal_out,
       calcuinter,
       ddsdata,
       ddsfqud,
       ddsreset,
       ddswclk,
       dumpoff,
       dumpon,
       interupt,
       k1,
       k2,
       pd_pulse_en,
       pulse_start,
       relay_close,
       relay_on,
       rt_sw,
       s_acq180,
       sd_acq_en,
       sigtimeup,
       soft_dump,
       sw_acq1,
       sw_acq2,
       syn_md_out,
       syn_md_tmp,
       xd
    );
input  [11:0] ADC;
input  OCX40MHz;
input  XRD;
input  ddsclkout;
input  gpio;
input  tri_ctrl;
input  [18:0] xa;
input  xwe;
input  zcs2;
output Acq_clk;
output GLA;
output Q1Q8;
output Q2Q7;
output Q3Q6;
output Q4Q5;
output cal_out;
output calcuinter;
output ddsdata;
output ddsfqud;
output ddsreset;
output ddswclk;
output dumpoff;
output dumpon;
output interupt;
output k1;
output k2;
output pd_pulse_en;
output pulse_start;
output [9:0] relay_close;
output [9:0] relay_on;
output rt_sw;
output s_acq180;
output sd_acq_en;
output sigtimeup;
output soft_dump;
output sw_acq1;
output sw_acq2;
output syn_md_out;
output syn_md_tmp;
inout  [15:0] xd;

    wire Signal_Noise_Acq_0_acq_clk, top_code_0_acqclken, net_27, 
        top_code_0_pluse_scale, scalestate_0_pluse_start, 
        plusestate_0_off_test, bri_dump_sw_0_off_test, 
        scalestate_0_off_test, bri_dump_sw_0_dump_start, 
        scalestate_0_dump_start, bri_dump_sw_0_phase_ctr, 
        scalestate_0_pn_out, top_code_0_pn_change, 
        bri_dump_sw_0_reset_out, net_45, top_code_0_pluse_rst, 
        bri_dump_sw_0_dumpoff_ctr, scalestate_0_dumpoff_ctr, 
        plusestate_0_tetw_pluse, bri_dump_sw_0_tetw_pluse, 
        bri_dump_sw_0_turn_delay, scalestate_0_ne_le, 
        top_code_0_bridge_load, \top_code_0_scaleddsdiv[0] , 
        \top_code_0_scaleddsdiv[1] , \top_code_0_scaleddsdiv[2] , 
        \top_code_0_scaleddsdiv[3] , \top_code_0_scaleddsdiv[4] , 
        \top_code_0_scaleddsdiv[5] , net_33, scanstate_0_calctrl, 
        top_code_0_cal_load, \top_code_0_cal_data[0] , 
        \top_code_0_cal_data[1] , \top_code_0_cal_data[2] , 
        \top_code_0_cal_data[3] , \top_code_0_cal_data[4] , 
        \top_code_0_cal_data[5] , top_code_0_sigrst, clock_10khz, 
        \top_code_0_sigtimedata[0] , \top_code_0_sigtimedata[1] , 
        \top_code_0_sigtimedata[2] , \top_code_0_sigtimedata[3] , 
        \top_code_0_sigtimedata[4] , \top_code_0_sigtimedata[5] , 
        \top_code_0_sigtimedata[6] , \top_code_0_sigtimedata[7] , 
        \top_code_0_sigtimedata[8] , \top_code_0_sigtimedata[9] , 
        \top_code_0_sigtimedata[10] , \top_code_0_sigtimedata[11] , 
        \top_code_0_sigtimedata[12] , \top_code_0_sigtimedata[13] , 
        \top_code_0_sigtimedata[14] , \top_code_0_sigtimedata[15] , 
        top_code_0_dds_load, top_code_0_dds_choice, 
        dds_change_0_dds_rst, dds_change_0_dds_conf, 
        \top_code_0_dds_configdata[0] , \top_code_0_dds_configdata[1] , 
        \top_code_0_dds_configdata[2] , \top_code_0_dds_configdata[3] , 
        \top_code_0_dds_configdata[4] , \top_code_0_dds_configdata[5] , 
        \top_code_0_dds_configdata[6] , \top_code_0_dds_configdata[7] , 
        \top_code_0_dds_configdata[8] , \top_code_0_dds_configdata[9] , 
        \top_code_0_dds_configdata[10] , 
        \top_code_0_dds_configdata[11] , 
        \top_code_0_dds_configdata[12] , 
        \top_code_0_dds_configdata[13] , 
        \top_code_0_dds_configdata[14] , 
        \top_code_0_dds_configdata[15] , \top_code_0_change[0] , 
        \top_code_0_change[1] , scalestate_0_dds_conf, 
        plusestate_0_dds_config, top_code_0_dump_sustain, net_40, 
        scalestate_0_dump_sustain_ctrl, 
        \top_code_0_dump_sustain_data[0] , 
        \top_code_0_dump_sustain_data[1] , 
        \top_code_0_dump_sustain_data[2] , 
        \top_code_0_dump_sustain_data[3] , state1ms_choice_0_reset_out, 
        state1ms_choice_0_dump_start, top_code_0_dumpload, 
        state1ms_choice_0_bri_cycle, bri_div_start_0, 
        \top_code_0_dump_cho_0[0] , \top_code_0_dump_cho_0[1] , 
        \top_code_0_dump_cho_0[2] , \top_code_0_dumpdata_0[0] , 
        \top_code_0_dumpdata_0[1] , \top_code_0_dumpdata_0[2] , 
        \top_code_0_dumpdata_0[3] , \top_code_0_dumpdata_0[4] , 
        \top_code_0_dumpdata_0[5] , \top_code_0_dumpdata_0[6] , 
        \top_code_0_dumpdata_0[7] , \top_code_0_dumpdata_0[8] , 
        \top_code_0_dumpdata_0[9] , \top_code_0_dumpdata_0[10] , 
        \top_code_0_dumpdata_0[11] , nsctrl_choice_0_dumponoff_rst, 
        nsctrl_choice_0_dumpoff_ctr, OR2_1_Y, OR2_2_Y, GPMI_0_code_en, 
        \Signal_Noise_Acq_0_dataout[12] , 
        \Signal_Noise_Acq_0_dataout[13] , 
        \Signal_Noise_Acq_0_dataout[14] , 
        \Signal_Noise_Acq_0_dataout[15] , top_code_0_pluse_noise_ctrl, 
        noisestate_0_n_acq, plusestate_0_pluse_acq, 
        n_acq_change_0_n_acq_start, top_code_0_noise_rst, 
        n_acq_change_0_n_rst_n, timer_top_0_clk_en_noise, 
        noisestate_0_dumpon_ctr, noisestate_0_dumpoff_ctr, 
        noisestate_0_soft_d, noisestate_0_rt_sw, noisestate_0_sw_acq2, 
        \noisestate_0_timecount[0] , \noisestate_0_timecount[1] , 
        \noisestate_0_timecount[2] , \noisestate_0_timecount[3] , 
        \noisestate_0_timecount[4] , \noisestate_0_timecount[5] , 
        \noisestate_0_timecount[6] , \noisestate_0_timecount[7] , 
        \noisestate_0_timecount[8] , \noisestate_0_timecount[9] , 
        \noisestate_0_timecount[10] , \noisestate_0_timecount[11] , 
        \noisestate_0_timecount[12] , \noisestate_0_timecount[13] , 
        \noisestate_0_timecount[14] , \noisestate_0_timecount[15] , 
        noisestate_0_state_over_n, top_code_0_nstateload, 
        top_code_0_nstatechoice, \top_code_0_noisedata[0] , 
        \top_code_0_noisedata[1] , \top_code_0_noisedata[2] , 
        \top_code_0_noisedata[3] , \top_code_0_noisedata[4] , 
        \top_code_0_noisedata[5] , \top_code_0_noisedata[6] , 
        \top_code_0_noisedata[7] , \top_code_0_noisedata[8] , 
        \top_code_0_noisedata[9] , \top_code_0_noisedata[10] , 
        \top_code_0_noisedata[11] , \top_code_0_noisedata[12] , 
        \top_code_0_noisedata[13] , \top_code_0_noisedata[14] , 
        \top_code_0_noisedata[15] , top_code_0_n_s_ctrl, 
        scanstate_0_soft_d, scanstate_0_rt_sw, scanstate_0_sw_acq2, 
        scanstate_0_state_over_n, scanstate_0_dds_conf, 
        scanstate_0_dumpoff_ctr, nsctrl_choice_0_soft_d, 
        nsctrl_choice_0_rt_sw, nsctrl_choice_0_sw_acq2, 
        nsctrl_choice_0_intertodsp, nsctrl_choice_0_dumpon_ctr, 
        top_code_0_pd_pluse_load, net_51, 
        \top_code_0_pd_pluse_choice[0] , 
        \top_code_0_pd_pluse_choice[1] , 
        \top_code_0_pd_pluse_choice[2] , 
        \top_code_0_pd_pluse_choice[3] , \top_code_0_pd_pluse_data[0] , 
        \top_code_0_pd_pluse_data[1] , \top_code_0_pd_pluse_data[2] , 
        \top_code_0_pd_pluse_data[3] , \top_code_0_pd_pluse_data[4] , 
        \top_code_0_pd_pluse_data[5] , \top_code_0_pd_pluse_data[6] , 
        \top_code_0_pd_pluse_data[7] , \top_code_0_pd_pluse_data[8] , 
        \top_code_0_pd_pluse_data[9] , \top_code_0_pd_pluse_data[10] , 
        \top_code_0_pd_pluse_data[11] , \top_code_0_pd_pluse_data[12] , 
        \top_code_0_pd_pluse_data[13] , \top_code_0_pd_pluse_data[14] , 
        \top_code_0_pd_pluse_data[15] , \top_code_0_bri_datain[0] , 
        \top_code_0_bri_datain[1] , \top_code_0_bri_datain[2] , 
        \top_code_0_bri_datain[3] , \top_code_0_bri_datain[4] , 
        \top_code_0_bri_datain[5] , \top_code_0_bri_datain[6] , 
        \top_code_0_bri_datain[7] , \top_code_0_bri_datain[8] , 
        \top_code_0_bri_datain[9] , \top_code_0_bri_datain[10] , 
        \top_code_0_bri_datain[11] , \top_code_0_bri_datain[12] , 
        \top_code_0_bri_datain[13] , \top_code_0_bri_datain[14] , 
        \top_code_0_bri_datain[15] , \top_code_0_halfdata_0[0] , 
        \top_code_0_halfdata_0[1] , \top_code_0_halfdata_0[2] , 
        \top_code_0_halfdata_0[3] , \top_code_0_halfdata_0[4] , 
        \top_code_0_halfdata_0[5] , \top_code_0_halfdata_0[6] , 
        \top_code_0_halfdata_0[7] , timer_top_0_clk_en_pluse, 
        plusestate_0_soft_d, plusestate_0_sw_acq1, 
        \plusestate_0_timecount[0] , \plusestate_0_timecount[1] , 
        \plusestate_0_timecount[2] , \plusestate_0_timecount[3] , 
        \plusestate_0_timecount[4] , \plusestate_0_timecount[5] , 
        \plusestate_0_timecount[6] , \plusestate_0_timecount[7] , 
        \plusestate_0_timecount[8] , \plusestate_0_timecount[9] , 
        \plusestate_0_timecount[10] , \plusestate_0_timecount[11] , 
        \plusestate_0_timecount[12] , \plusestate_0_timecount[13] , 
        \plusestate_0_timecount[14] , \plusestate_0_timecount[15] , 
        \top_code_0_plusedata[0] , \top_code_0_plusedata[1] , 
        \top_code_0_plusedata[2] , \top_code_0_plusedata[3] , 
        \top_code_0_plusedata[4] , \top_code_0_plusedata[5] , 
        \top_code_0_plusedata[6] , \top_code_0_plusedata[7] , 
        \top_code_0_plusedata[8] , \top_code_0_plusedata[9] , 
        \top_code_0_plusedata[10] , \top_code_0_plusedata[11] , 
        \top_code_0_plusedata[12] , \top_code_0_plusedata[13] , 
        \top_code_0_plusedata[14] , \top_code_0_plusedata[15] , 
        top_code_0_pluseload, top_code_0_pluse_lc, 
        plusestate_0_state_over_n, s_acq_change_0_s_load, 
        top_code_0_s_load, scalestate_0_load_out, s_acq_change_0_s_rst, 
        \s_acq_change_0_s_acqnum[0] , \s_acq_change_0_s_acqnum[1] , 
        \s_acq_change_0_s_acqnum[2] , \s_acq_change_0_s_acqnum[3] , 
        \s_acq_change_0_s_acqnum[4] , \s_acq_change_0_s_acqnum[5] , 
        \s_acq_change_0_s_acqnum[6] , \s_acq_change_0_s_acqnum[7] , 
        \s_acq_change_0_s_acqnum[8] , \s_acq_change_0_s_acqnum[9] , 
        \s_acq_change_0_s_acqnum[10] , \s_acq_change_0_s_acqnum[11] , 
        \s_acq_change_0_s_acqnum[12] , \s_acq_change_0_s_acqnum[13] , 
        \s_acq_change_0_s_acqnum[14] , \s_acq_change_0_s_acqnum[15] , 
        \top_code_0_s_acqnum_2[0] , \top_code_0_s_acqnum_2[1] , 
        \top_code_0_s_acqnum_2[2] , \top_code_0_s_acqnum_2[3] , 
        \top_code_0_s_acqnum_2[4] , \top_code_0_s_acqnum_2[5] , 
        \top_code_0_s_acqnum_2[6] , \top_code_0_s_acqnum_2[7] , 
        \top_code_0_s_acqnum_2[8] , \top_code_0_s_acqnum_2[9] , 
        \top_code_0_s_acqnum_2[10] , \top_code_0_s_acqnum_2[11] , 
        \top_code_0_s_acqnum_2[12] , \top_code_0_s_acqnum_2[13] , 
        \top_code_0_s_acqnum_2[14] , \top_code_0_s_acqnum_2[15] , 
        \scalestate_0_s_acqnum[0] , \scalestate_0_s_acqnum[1] , 
        \scalestate_0_s_acqnum[2] , \scalestate_0_s_acqnum[3] , 
        \scalestate_0_s_acqnum[4] , \scalestate_0_s_acqnum[5] , 
        \scalestate_0_s_acqnum[6] , \scalestate_0_s_acqnum[7] , 
        \scalestate_0_s_acqnum[8] , \scalestate_0_s_acqnum[9] , 
        \scalestate_0_s_acqnum[10] , \scalestate_0_s_acqnum[11] , 
        \s_acq_change_0_s_stripnum[0] , \s_acq_change_0_s_stripnum[1] , 
        \s_acq_change_0_s_stripnum[2] , \s_acq_change_0_s_stripnum[3] , 
        \s_acq_change_0_s_stripnum[4] , \s_acq_change_0_s_stripnum[5] , 
        \s_acq_change_0_s_stripnum[6] , \s_acq_change_0_s_stripnum[7] , 
        \s_acq_change_0_s_stripnum[8] , \s_acq_change_0_s_stripnum[9] , 
        \s_acq_change_0_s_stripnum[10] , 
        \s_acq_change_0_s_stripnum[11] , \scalestate_0_strippluse[0] , 
        \scalestate_0_strippluse[1] , \scalestate_0_strippluse[2] , 
        \scalestate_0_strippluse[3] , \scalestate_0_strippluse[4] , 
        \scalestate_0_strippluse[5] , \scalestate_0_strippluse[6] , 
        \scalestate_0_strippluse[7] , \scalestate_0_strippluse[8] , 
        \scalestate_0_strippluse[9] , \scalestate_0_strippluse[10] , 
        \scalestate_0_strippluse[11] , timer_top_0_clk_en_scale, 
        top_code_0_scale_rst, scalestate_0_soft_d, scalestate_0_rt_sw, 
        scalestate_0_sw_acq1, scalestate_0_sw_acq2, 
        \scalestate_0_timecount[0] , \scalestate_0_timecount[1] , 
        \scalestate_0_timecount[2] , \scalestate_0_timecount[3] , 
        \scalestate_0_timecount[4] , \scalestate_0_timecount[5] , 
        \scalestate_0_timecount[7] , \scalestate_0_timecount[8] , 
        \scalestate_0_timecount[9] , \scalestate_0_timecount[10] , 
        \scalestate_0_timecount[11] , \scalestate_0_timecount[12] , 
        \scalestate_0_timecount[13] , \scalestate_0_timecount[14] , 
        \scalestate_0_timecount[15] , \scalestate_0_timecount[16] , 
        \scalestate_0_timecount[17] , \scalestate_0_timecount[18] , 
        \scalestate_0_timecount[19] , \scalestate_0_timecount[20] , 
        \scalestate_0_timecount[21] , scalestate_0_s_acq, 
        \top_code_0_scaledatain[0] , \top_code_0_scaledatain[1] , 
        \top_code_0_scaledatain[2] , \top_code_0_scaledatain[3] , 
        \top_code_0_scaledatain[4] , \top_code_0_scaledatain[5] , 
        \top_code_0_scaledatain[6] , \top_code_0_scaledatain[7] , 
        \top_code_0_scaledatain[8] , \top_code_0_scaledatain[9] , 
        \top_code_0_scaledatain[10] , \top_code_0_scaledatain[11] , 
        \top_code_0_scaledatain[12] , \top_code_0_scaledatain[13] , 
        \top_code_0_scaledatain[14] , \top_code_0_scaledatain[15] , 
        top_code_0_scaleload, \top_code_0_scalechoice_0[0] , 
        \top_code_0_scalechoice_0[1] , \top_code_0_scalechoice_0[2] , 
        \top_code_0_scalechoice_0[3] , \top_code_0_scalechoice_0[4] , 
        top_code_0_inv_turn, scalestate_0_tetw_pluse, 
        scalestate_0_long_opentime, scan_scale_sw_0_s_start, 
        scanstate_0_s_acq, timer_top_0_clk_en_scan, 
        \scanstate_0_timecount[0] , \scanstate_0_timecount[1] , 
        \scanstate_0_timecount[2] , \scanstate_0_timecount[3] , 
        \scanstate_0_timecount[4] , \scanstate_0_timecount[5] , 
        \scanstate_0_timecount[6] , \scanstate_0_timecount[7] , 
        \scanstate_0_timecount[8] , \scanstate_0_timecount[9] , 
        \scanstate_0_timecount[10] , \scanstate_0_timecount[11] , 
        \scanstate_0_timecount[12] , \scanstate_0_timecount[13] , 
        \scanstate_0_timecount[14] , \scanstate_0_timecount[15] , 
        top_code_0_scanload, \top_code_0_scandata[0] , 
        \top_code_0_scandata[1] , \top_code_0_scandata[2] , 
        \top_code_0_scandata[3] , \top_code_0_scandata[4] , 
        \top_code_0_scandata[5] , \top_code_0_scandata[6] , 
        \top_code_0_scandata[7] , \top_code_0_scandata[8] , 
        \top_code_0_scandata[9] , \top_code_0_scandata[10] , 
        \top_code_0_scandata[11] , \top_code_0_scandata[12] , 
        \top_code_0_scandata[13] , \top_code_0_scandata[14] , 
        \top_code_0_scandata[15] , top_code_0_scanchoice, 
        top_code_0_sd_sacq_load, \top_code_0_sd_sacq_choice[0] , 
        \top_code_0_sd_sacq_choice[1] , \top_code_0_sd_sacq_choice[2] , 
        \top_code_0_sd_sacq_choice[3] , \top_code_0_sd_sacq_data[0] , 
        \top_code_0_sd_sacq_data[1] , \top_code_0_sd_sacq_data[2] , 
        \top_code_0_sd_sacq_data[3] , \top_code_0_sd_sacq_data[4] , 
        \top_code_0_sd_sacq_data[5] , \top_code_0_sd_sacq_data[6] , 
        \top_code_0_sd_sacq_data[7] , \top_code_0_sd_sacq_data[8] , 
        \top_code_0_sd_sacq_data[9] , \top_code_0_sd_sacq_data[10] , 
        \top_code_0_sd_sacq_data[11] , \top_code_0_sd_sacq_data[12] , 
        \top_code_0_sd_sacq_data[13] , \top_code_0_sd_sacq_data[14] , 
        \top_code_0_sd_sacq_data[15] , top_code_0_n_load, 
        top_code_0_RAM_Rd_rst, top_code_0_n_rd_en, 
        \top_code_0_n_acqnum_2[0] , \top_code_0_n_acqnum_2[1] , 
        \top_code_0_n_acqnum_2[2] , \top_code_0_n_acqnum_2[3] , 
        \top_code_0_n_acqnum_2[4] , \top_code_0_n_acqnum_2[5] , 
        \top_code_0_n_acqnum_2[6] , \top_code_0_n_acqnum_2[7] , 
        \top_code_0_n_acqnum_2[8] , \top_code_0_n_acqnum_2[9] , 
        \top_code_0_n_acqnum_2[10] , \top_code_0_n_acqnum_2[11] , 
        \top_code_0_n_divnum_0[0] , \top_code_0_n_divnum_0[1] , 
        \top_code_0_n_divnum_0[2] , \top_code_0_n_divnum_0[3] , 
        \top_code_0_n_divnum_0[4] , \top_code_0_n_divnum_0[5] , 
        \top_code_0_n_divnum_0[6] , \top_code_0_n_divnum_0[7] , 
        \top_code_0_n_divnum_0[8] , \top_code_0_n_divnum_0[9] , 
        \top_code_0_s_periodnum[0] , \top_code_0_s_periodnum[1] , 
        \top_code_0_s_periodnum[2] , \top_code_0_s_periodnum[3] , 
        \top_code_0_s_addchoice[0] , \top_code_0_s_addchoice[1] , 
        \top_code_0_s_addchoice[2] , \top_code_0_s_addchoice[3] , 
        \top_code_0_s_addchoice[4] , top_code_0_state_1ms_start, 
        state_1ms_0_pluse_start, state_1ms_0_dump_start, 
        state_1ms_0_reset_out, state_1ms_0_bri_cycle, 
        state_1ms_0_rt_sw, rt_sw_net_0, state_1ms_0_soft_dump, 
        soft_dump_net_0, timer_top_0_clk_en_st1ms, 
        top_code_0_state_1ms_rst_n, top_code_0_state_1ms_load, 
        \top_code_0_state_1ms_lc[0] , \top_code_0_state_1ms_lc[1] , 
        \top_code_0_state_1ms_lc[2] , \top_code_0_state_1ms_lc[3] , 
        \top_code_0_state_1ms_data[0] , \top_code_0_state_1ms_data[1] , 
        \top_code_0_state_1ms_data[2] , \top_code_0_state_1ms_data[3] , 
        \top_code_0_state_1ms_data[4] , \top_code_0_state_1ms_data[5] , 
        \top_code_0_state_1ms_data[6] , \top_code_0_state_1ms_data[7] , 
        \top_code_0_state_1ms_data[8] , \top_code_0_state_1ms_data[9] , 
        \top_code_0_state_1ms_data[10] , 
        \top_code_0_state_1ms_data[11] , 
        \top_code_0_state_1ms_data[12] , 
        \top_code_0_state_1ms_data[13] , 
        \top_code_0_state_1ms_data[14] , 
        \top_code_0_state_1ms_data[15] , \state_1ms_0_timecount[0] , 
        \state_1ms_0_timecount[1] , \state_1ms_0_timecount[2] , 
        \state_1ms_0_timecount[3] , \state_1ms_0_timecount[4] , 
        \state_1ms_0_timecount[5] , \state_1ms_0_timecount[6] , 
        \state_1ms_0_timecount[7] , \state_1ms_0_timecount[8] , 
        \state_1ms_0_timecount[9] , \state_1ms_0_timecount[10] , 
        \state_1ms_0_timecount[11] , \state_1ms_0_timecount[12] , 
        \state_1ms_0_timecount[13] , \state_1ms_0_timecount[14] , 
        \state_1ms_0_timecount[15] , \state_1ms_0_timecount[16] , 
        \state_1ms_0_timecount[17] , \state_1ms_0_timecount[18] , 
        \state_1ms_0_timecount[19] , top_code_0_scale_start, 
        top_code_0_scan_start, top_code_0_noise_start, 
        top_code_0_pluse_str, \GPMI_0.tri_state_0.xd_1 , 
        \Signal_Noise_Acq_0_dataout[0] , 
        \Signal_Noise_Acq_0_dataout[1] , 
        \Signal_Noise_Acq_0_dataout[2] , 
        \Signal_Noise_Acq_0_dataout[3] , 
        \Signal_Noise_Acq_0_dataout[4] , 
        \Signal_Noise_Acq_0_dataout[5] , 
        \Signal_Noise_Acq_0_dataout[6] , 
        \Signal_Noise_Acq_0_dataout[7] , 
        \Signal_Noise_Acq_0_dataout[8] , 
        \Signal_Noise_Acq_0_dataout[9] , 
        \Signal_Noise_Acq_0_dataout[10] , 
        \Signal_Noise_Acq_0_dataout[11] , \i_0_0[1] , \i_6[1] , 
        DUMP_ON_0_dump_on, DUMP_OFF_1_dump_off, DUMP_OFF_0_dump_off, 
        DUMP_0_dump_off, DUMP_0_dump_on, \xd_in[0] , \xd_in[1] , 
        \xd_in[2] , \xd_in[3] , \xd_in[4] , \xd_in[5] , \xd_in[6] , 
        \xd_in[7] , \xd_in[8] , \xd_in[9] , \xd_in[10] , \xd_in[11] , 
        \xd_in[12] , \xd_in[13] , \xd_in[14] , \xd_in[15] , \ADC_c[0] , 
        \ADC_c[1] , \ADC_c[2] , \ADC_c[3] , \ADC_c[4] , \ADC_c[5] , 
        \ADC_c[6] , \ADC_c[7] , \ADC_c[8] , \ADC_c[9] , \ADC_c[10] , 
        \ADC_c[11] , XRD_c, ddsclkout_c, gpio_c, tri_ctrl_c, \xa_c[0] , 
        \xa_c[1] , \xa_c[2] , \xa_c[3] , \xa_c[4] , \xa_c[5] , 
        \xa_c[6] , \xa_c[7] , \xa_c[8] , \xa_c[9] , \xa_c[10] , 
        \xa_c[11] , \xa_c[12] , \xa_c[13] , \xa_c[14] , \xa_c[15] , 
        \xa_c[16] , \xa_c[17] , \xa_c[18] , xwe_c, zcs2_c, Acq_clk_c, 
        GLA_net_1, Q3Q6_c, Q4Q5_c, cal_out_c, calcuinter_c, dumpoff_c, 
        dumpon_c, interupt_c, k1_c, k2_c, pd_pulse_en_c, pulse_start_c, 
        \relay_close_c[0] , \relay_close_c[1] , \relay_close_c[2] , 
        \relay_close_c[3] , \relay_close_c[4] , \relay_close_c[5] , 
        \relay_close_c[6] , \relay_close_c[7] , \relay_close_c[8] , 
        \relay_close_c[9] , \relay_on_c[0] , \relay_on_c[1] , 
        \relay_on_c[2] , \relay_on_c[3] , \relay_on_c[4] , 
        \relay_on_c[5] , \relay_on_c[6] , \relay_on_c[7] , 
        \relay_on_c[8] , \relay_on_c[9] , s_acq180_c, sd_acq_en_c, 
        sigtimeup_c, sw_acq1_c, sw_acq2_c, syn_md_out_c, syn_md_tmp_c, 
        \GPMI_0_dataout[0] , \GPMI_0_dataout[1] , \GPMI_0_dataout[2] , 
        \GPMI_0_dataout[3] , \GPMI_0_dataout[4] , \GPMI_0_dataout[5] , 
        \GPMI_0_dataout[6] , \GPMI_0_dataout[7] , PLUSE_0_bri_cycle, 
        \dds_change_0.un1_change_2 , \GPMI_0_dataout[11] , 
        \GPMI_0_dataout[8] , \GPMI_0_dataout[9] , \GPMI_0_dataout[10] , 
        \GPMI_0_dataout[12] , \GPMI_0_dataout[13] , 
        \GPMI_0_dataout[14] , \GPMI_0_dataout[15] , clk_4f_en, 
        clk_4f_en_0, \GPMI_0_dataout_0[3] , \GPMI_0_dataout_0[2] , 
        \GPMI_0_dataout_0[1] , \GPMI_0_dataout_0[0] , 
        top_code_0_state_1ms_rst_n_0, \top_code_0_s_addchoice_0[4] , 
        \top_code_0_s_addchoice_1[4] , \top_code_0_s_addchoice_2[4] , 
        \top_code_0_s_addchoice_3[4] , \top_code_0_s_addchoice_4[4] , 
        \top_code_0_s_addchoice_5[4] , \top_code_0_s_addchoice_0[2] , 
        \top_code_0_s_addchoice_0[1] , \top_code_0_s_addchoice_1[1] , 
        \top_code_0_s_addchoice_0[0] , \top_code_0_s_addchoice_1[0] , 
        \top_code_0_s_addchoice_2[0] , \top_code_0_s_addchoice_3[0] , 
        \top_code_0_s_addchoice_4[0] , \top_code_0_scalechoice_0_0[0] , 
        \top_code_0_scaledatain_0[3] , \top_code_0_scaledatain_0[2] , 
        \top_code_0_scaledatain_0[1] , \top_code_0_scaledatain_0[0] , 
        top_code_0_scale_rst_0, top_code_0_scale_rst_1, 
        top_code_0_scale_rst_2, top_code_0_scale_rst_3, 
        top_code_0_scale_rst_4, top_code_0_scale_rst_5, 
        timer_top_0_clk_en_scale_0, s_acq_change_0_s_load_0, 
        top_code_0_n_s_ctrl_0, top_code_0_n_s_ctrl_1, 
        n_acq_change_0_n_rst_n_0, top_code_0_noise_rst_0, 
        \top_code_0_change_0[1] , \top_code_0_change_0[0] , net_33_0, 
        top_code_0_bridge_load_0, top_code_0_pluse_rst_0, 
        bri_dump_sw_0_reset_out_0, \GPMI_0_dataout_0[4] , 
        \state1ms_choice_0/bri_cycle_RNO_net_1 , 
        \state1ms_choice_0/bri_cycle_5 , 
        \state1ms_choice_0/dump_start_RNO_1 , 
        \state1ms_choice_0/dump_start_5 , 
        \state1ms_choice_0/pluse_start_RNO_1 , 
        \state1ms_choice_0/pluse_start_5 , 
        \state1ms_choice_0/reset_out_RNO_0_net_1 , 
        \state1ms_choice_0/reset_out_5 , 
        \state1ms_choice_0/soft_dump_4 , \state1ms_choice_0/rt_sw_4 , 
        \top_code_0/pluse_rst_0_0_RNIO7ND3_net_1 , \top_code_0/N_62 , 
        \top_code_0/scan_rst_RNIMNCI3_net_1 , 
        \top_code_0/change_1_sqmuxa , 
        \top_code_0/noise_rst_0_0_RNIDOO43_net_1 , \top_code_0/N_76 , 
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 , 
        \top_code_0/scaledatain_1_sqmuxa , 
        \top_code_0/scalechoice_1_sqmuxa , 
        \top_code_0/s_addchoice_1_sqmuxa , 
        \top_code_0/state_1ms_rst_n_0_0_RNI848T5_net_1 , 
        \top_code_0/N_112_reto , \top_code_0/N_112 , 
        \top_code_0/un1_xa_4_reto , \top_code_0/un1_xa_4 , 
        \top_code_0/top_code_0_state_1ms_start_reto , 
        \top_code_0/N_795_reto , \top_code_0/N_110_reto , 
        \top_code_0/N_110 , \top_code_0/xa_c_reto[0] , 
        \top_code_0/top_code_0_scale_start_reto , 
        \top_code_0/N_797_reto , \top_code_0/N_114_reto , 
        \top_code_0/N_114 , \top_code_0/un1_xa_13_reto , 
        \top_code_0/un1_xa_13 , 
        \top_code_0/top_code_0_noise_start_reto , 
        \top_code_0/N_799_reto , \top_code_0/N_108_reto , 
        \top_code_0/N_108 , \top_code_0/un1_xa_10_reto , 
        \top_code_0/un1_xa_10 , 
        \top_code_0/top_code_0_scan_start_reto , 
        \top_code_0/N_796_reto , \top_code_0/net_27_reto , 
        \top_code_0/N_327 , \top_code_0/N_171 , 
        \top_code_0/un1_state_1ms_rst_n117_44_i_a2_0 , 
        \top_code_0/N_162 , \top_code_0/N_174 , \top_code_0/N_329 , 
        \top_code_0/un1_state_1ms_rst_n117_47_i_a2_0 , 
        \top_code_0/N_328 , \top_code_0/N_330 , \top_code_0/N_137 , 
        \top_code_0/un1_xa_30_0_o2_0_net_1 , \top_code_0/N_139 , 
        \top_code_0/N_192 , \top_code_0/N_334 , 
        \top_code_0/scandata_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_157 , 
        \top_code_0/noisedata_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_333 , 
        \top_code_0/state_1ms_data_1_sqmuxa_0_a2_1_net_1 , 
        \top_code_0/n_acqnum_1_sqmuxa_0_a2_0 , \top_code_0/N_154 , 
        \top_code_0/N_147 , \top_code_0/N_163 , 
        \top_code_0/plusedata_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_340 , 
        \top_code_0/s_addchoice_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_144 , \top_code_0/N_164 , 
        \top_code_0/state_1ms_lc_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/s_periodnum_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_159 , \top_code_0/N_150 , \top_code_0/N_165 , 
        \top_code_0/N_161 , \top_code_0/N_332 , \top_code_0/N_149 , 
        \top_code_0/un1_state_1ms_rst_n117_i_a2_0_net_1 , 
        \top_code_0/relay_close_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/N_337 , 
        \top_code_0/relay_on_1_sqmuxa_0_a2_0_net_1 , 
        \top_code_0/un1_state_1ms_rst_n117_43_i_a3_0_0_net_1 , 
        \top_code_0/N_140 , 
        \top_code_0/un1_state_1ms_rst_n117_18_i_o2_0_net_1 , 
        \top_code_0/un1_state_1ms_rst_n117_43_i_a2_1_1_net_1 , 
        \top_code_0/un1_state_1ms_rst_n117_43_i_a2_0_0_net_1 , 
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_3_net_1 , 
        \top_code_0/N_13 , 
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_1 , 
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_2 , 
        \top_code_0/N_127 , 
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_4 , 
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_2 , 
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_3 , 
        \top_code_0/N_158 , 
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_5_net_1 , 
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_3_net_1 , 
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_4_net_1 , 
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_1_net_1 , 
        \top_code_0/un1_xa_4_0_a2_1 , \top_code_0/un1_xa_49_0_a2_1 , 
        \top_code_0/relay_on_1_sqmuxa , 
        \top_code_0/state_1ms_data_1_sqmuxa , \top_code_0/N_152 , 
        \top_code_0/state_1ms_lc_1_sqmuxa , \top_code_0/N_326 , 
        \top_code_0/N_325 , \top_code_0/N_320 , \top_code_0/N_169 , 
        \top_code_0/sd_sacq_choice_1_sqmuxa , \top_code_0/N_331 , 
        \top_code_0/N_336 , \top_code_0/plusedata_1_sqmuxa , 
        \top_code_0/n_acqnum_1_sqmuxa , \top_code_0/un1_xa_49 , 
        \top_code_0/N_339 , \top_code_0/N_11 , \top_code_0/N_11_3 , 
        \top_code_0/N_12 , \top_code_0/N_167 , \top_code_0/N_321 , 
        \top_code_0/N_148 , \top_code_0/N_302 , \top_code_0/N_258 , 
        \top_code_0/N_259 , \top_code_0/N_264 , 
        \top_code_0/sd_sacq_data_1_sqmuxa , 
        \top_code_0/scandata_1_sqmuxa , \top_code_0/N_151 , 
        \top_code_0/N_142 , \top_code_0/s_periodnum_1_sqmuxa , 
        \top_code_0/noisedata_1_sqmuxa , \top_code_0/un1_xa_10_2 , 
        \top_code_0/relay_close_1_sqmuxa , \top_code_0/N_802 , 
        \top_code_0/N_122 , \top_code_0/N_808 , \top_code_0/N_262 , 
        \top_code_0/dump_sustain_RNO_net_1 , 
        \top_code_0/inv_turn_RNO_net_1 , 
        \top_code_0/relay_close_RNO[0]_net_1 , \top_code_0/N_819 , 
        \top_code_0/relay_close_RNO[1]_net_1 , \top_code_0/N_820 , 
        \top_code_0/relay_close_RNO[2]_net_1 , \top_code_0/N_821 , 
        \top_code_0/relay_close_RNO[3]_net_1 , \top_code_0/N_822 , 
        \top_code_0/relay_close_RNO[4]_net_1 , \top_code_0/N_823 , 
        \top_code_0/relay_close_RNO[5]_net_1 , \top_code_0/N_824 , 
        \top_code_0/relay_close_RNO[6]_net_1 , \top_code_0/N_825 , 
        \top_code_0/relay_close_RNO[7]_net_1 , \top_code_0/N_826 , 
        \top_code_0/relay_close_RNO[8]_net_1 , \top_code_0/N_827 , 
        \top_code_0/relay_close_RNO[9]_net_1 , \top_code_0/N_828 , 
        \top_code_0/relay_on_RNO[0]_net_1 , \top_code_0/N_809 , 
        \top_code_0/relay_on_RNO[1]_net_1 , \top_code_0/N_810 , 
        \top_code_0/relay_on_RNO[2]_net_1 , \top_code_0/N_811 , 
        \top_code_0/relay_on_RNO[3]_net_1 , \top_code_0/N_812 , 
        \top_code_0/relay_on_RNO[4]_net_1 , \top_code_0/N_813 , 
        \top_code_0/relay_on_RNO[5]_net_1 , \top_code_0/N_814 , 
        \top_code_0/relay_on_RNO[6]_net_1 , \top_code_0/N_815 , 
        \top_code_0/relay_on_RNO[7]_net_1 , \top_code_0/N_816 , 
        \top_code_0/relay_on_RNO[8]_net_1 , \top_code_0/N_817 , 
        \top_code_0/relay_on_RNO[9]_net_1 , \top_code_0/N_818 , 
        \top_code_0/N_219 , \top_code_0/N_160 , \top_code_0/N_218 , 
        \top_code_0/N_217 , \top_code_0/N_207 , \top_code_0/N_155 , 
        \top_code_0/N_203 , \top_code_0/N_202 , \top_code_0/N_199 , 
        \top_code_0/N_197 , \top_code_0/N_322 , \top_code_0/N_106 , 
        \top_code_0/N_314 , \top_code_0/N_100 , \top_code_0/N_308 , 
        \top_code_0/N_96 , \top_code_0/N_304 , \top_code_0/N_92 , 
        \top_code_0/N_300 , \top_code_0/N_90 , \top_code_0/N_175 , 
        \top_code_0/N_297 , \top_code_0/N_86 , \top_code_0/N_176 , 
        \top_code_0/N_293 , \top_code_0/N_84 , \top_code_0/N_291 , 
        \top_code_0/N_82 , \top_code_0/N_290 , \top_code_0/N_70 , 
        \top_code_0/N_278 , \top_code_0/N_60 , \top_code_0/N_268 , 
        \top_code_0/n_divnum_1_sqmuxa , \top_code_0/dumpdata_1_sqmuxa , 
        \top_code_0/dump_cho_1_sqmuxa , 
        \top_code_0/bri_datain_1_sqmuxa , 
        \top_code_0/pd_pluse_choice_1_sqmuxa , 
        \top_code_0/sigtimedata_1_sqmuxa_1 , 
        \top_code_0/pd_pluse_data_1_sqmuxa , 
        \top_code_0/dds_configdata_1_sqmuxa_1 , \top_code_0/N_266 , 
        \top_code_0/N_274 , \top_code_0/N_58 , \top_code_0/N_206 , 
        \top_code_0/N_66 , \top_code_0/N_205 , \top_code_0/N_284 , 
        \top_code_0/s_acqnum_1_sqmuxa_1 , \top_code_0/N_198 , 
        \top_code_0/dds_configdata_1_sqmuxa , \top_code_0/N_276 , 
        \top_code_0/N_286 , \top_code_0/N_288 , \top_code_0/N_319 , 
        \top_code_0/N_190 , \top_code_0/N_68 , \top_code_0/N_200 , 
        \top_code_0/N_78 , \top_code_0/N_210 , \top_code_0/N_80 , 
        \top_code_0/N_211 , \top_code_0/N_803 , \top_code_0/N_804 , 
        \top_code_0/N_805 , \top_code_0/N_280 , \top_code_0/N_72 , 
        \top_code_0/N_201 , \top_code_0/N_94 , \top_code_0/N_196 , 
        \top_code_0/N_801 , \top_code_0/k2_RNO_net_1 , 
        \top_code_0/N_806 , \top_code_0/k1_RNO_net_1 , 
        \top_code_0/N_807 , \top_code_0/N_295 , \top_code_0/N_88 , 
        \top_code_0/N_798 , \top_code_0/N_116 , 
        \top_code_0/pluse_str_RNO_net_1 , \top_code_0/N_208 , 
        \top_code_0/N_98 , \top_code_0/N_306 , 
        \top_code_0/sigtimedata_1_sqmuxa , 
        \top_code_0/s_acqnum_1_sqmuxa , 
        \top_code_0/dump_sustain_data_1_sqmuxa , 
        \top_code_0/cal_data_1_sqmuxa_1 , \top_code_0/N_312 , 
        \top_code_0/N_104 , \top_code_0/N_209 , \top_code_0/N_310 , 
        \top_code_0/N_102 , \top_code_0/N_195 , \top_code_0/N_800 , 
        \top_code_0/un1_xa_2 , \top_code_0/cal_data_1_sqmuxa , 
        \top_code_0/halfdata_1_sqmuxa , 
        \top_code_0/scaleddsdiv_1_sqmuxa , \top_code_0/N_270 , 
        \top_code_0/N_272 , \top_code_0/N_282 , \top_code_0/N_216 , 
        \top_code_0/N_64 , \top_code_0/N_204 , \top_code_0/N_74 , 
        \scan_scale_sw_0/s_start_RNO_net_1 , \scan_scale_sw_0/N_26 , 
        \scan_scale_sw_0/s_start_5 , \DDS_0/count[0] , 
        \DDS_0/count[1] , \DDS_0/count[2] , \DDS_0/count[3] , 
        \DDS_0/count[4] , \DDS_0/count[5] , \DDS_0/count[6] , 
        \DDS_0/count[7] , \DDS_0/dds_state_0_state_over , \DDS_0/i[0] , 
        \DDS_0/i[1] , \DDS_0/i[2] , \DDS_0/i[3] , 
        \DDS_0/dds_timer_0/count_15_0 , 
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 , 
        \DDS_0/dds_timer_0/N_36 , \DDS_0/dds_timer_0/count_c4 , 
        \DDS_0/dds_timer_0/count_n2 , \DDS_0/dds_timer_0/count_c1 , 
        \DDS_0/dds_timer_0/count_n3 , \DDS_0/dds_timer_0/count_c2 , 
        \DDS_0/dds_timer_0/count_n4 , \DDS_0/dds_timer_0/count_c3 , 
        \DDS_0/dds_timer_0/count_n5 , \DDS_0/dds_timer_0/count_n6 , 
        \DDS_0/dds_timer_0/count_n6_tz , \DDS_0/dds_timer_0/count_n0 , 
        \DDS_0/dds_timer_0/count_n1 , \DDS_0/dds_timer_0/count_n7 , 
        \DDS_0/dds_state_0/N_569_1 , \DDS_0/dds_state_0/N_569_0 , 
        \DDS_0/dds_state_0/N_538_1 , \DDS_0/dds_state_0/N_538_0 , 
        \DDS_0/dds_state_0/N_535_0 , \DDS_0/dds_state_0/N_534_0 , 
        \DDS_0/dds_state_0/para_1_sqmuxa_1_0 , 
        \DDS_0/dds_state_0/w_clk_reg_net_1 , 
        \DDS_0/dds_state_0/para_9_i_1[16] , 
        \DDS_0/dds_state_0/para[16]_net_1 , \DDS_0/dds_state_0/N_294 , 
        \DDS_0/dds_state_0/para_9_i_1[13] , 
        \DDS_0/dds_state_0/para[13]_net_1 , \DDS_0/dds_state_0/N_334 , 
        \DDS_0/dds_state_0/para_9_i_1[29] , \DDS_0/dds_state_0/N_569 , 
        \DDS_0/dds_state_0/N_482 , \DDS_0/dds_state_0/para_9_i_1[24] , 
        \DDS_0/dds_state_0/N_303 , \DDS_0/dds_state_0/para_9_i_1[26] , 
        \DDS_0/dds_state_0/N_470 , \DDS_0/dds_state_0/para_9_i_1[30] , 
        \DDS_0/dds_state_0/N_514 , \DDS_0/dds_state_0/para_9_i_1[23] , 
        \DDS_0/dds_state_0/N_299 , \DDS_0/dds_state_0/para_9_i_1[11] , 
        \DDS_0/dds_state_0/para[11]_net_1 , \DDS_0/dds_state_0/N_325 , 
        \DDS_0/dds_state_0/para_9_i_0[31] , 
        \DDS_0/dds_state_0/para_reg[31]_net_1 , 
        \DDS_0/dds_state_0/N_520 , \DDS_0/dds_state_0/para_9_i_1[2] , 
        \DDS_0/dds_state_0/para[2]_net_1 , \DDS_0/dds_state_0/N_485 , 
        \DDS_0/dds_state_0/para_9_i_1[14] , 
        \DDS_0/dds_state_0/para[14]_net_1 , \DDS_0/dds_state_0/N_461 , 
        \DDS_0/dds_state_0/para_9_i_1[32] , \DDS_0/dds_state_0/N_312 , 
        \DDS_0/dds_state_0/para_9_i_1[20] , \DDS_0/dds_state_0/N_466 , 
        \DDS_0/dds_state_0/para_9_i_1[27] , \DDS_0/dds_state_0/N_474 , 
        \DDS_0/dds_state_0/para_9_i_1[19] , \DDS_0/dds_state_0/N_506 , 
        \DDS_0/dds_state_0/para_9_i_0_1[6] , 
        \DDS_0/dds_state_0/para[6]_net_1 , \DDS_0/dds_state_0/N_274 , 
        \DDS_0/dds_state_0/para_9_i_1[28] , \DDS_0/dds_state_0/N_478 , 
        \DDS_0/dds_state_0/para_9_i_0_1[1] , 
        \DDS_0/dds_state_0/para[1]_net_1 , \DDS_0/dds_state_0/N_278 , 
        \DDS_0/dds_state_0/para_9_i_1[15] , 
        \DDS_0/dds_state_0/para[15]_net_1 , \DDS_0/dds_state_0/N_493 , 
        \DDS_0/dds_state_0/para_9_i_1[25] , \DDS_0/dds_state_0/N_307 , 
        \DDS_0/dds_state_0/para_9_i_1[12] , 
        \DDS_0/dds_state_0/para[12]_net_1 , \DDS_0/dds_state_0/N_329 , 
        \DDS_0/dds_state_0/para_9_i_1[10] , 
        \DDS_0/dds_state_0/para[10]_net_1 , \DDS_0/dds_state_0/N_290 , 
        \DDS_0/dds_state_0/para_9_i_1[3] , 
        \DDS_0/dds_state_0/para[3]_net_1 , \DDS_0/dds_state_0/N_489 , 
        \DDS_0/dds_state_0/para_9_i_1[18] , \DDS_0/dds_state_0/N_502 , 
        \DDS_0/dds_state_0/para_9_i_1[4] , 
        \DDS_0/dds_state_0/para[4]_net_1 , \DDS_0/dds_state_0/N_315 , 
        \DDS_0/dds_state_0/para_9_i_1[9] , 
        \DDS_0/dds_state_0/para[9]_net_1 , \DDS_0/dds_state_0/N_286 , 
        \DDS_0/dds_state_0/para_9_i_1[8] , 
        \DDS_0/dds_state_0/para[8]_net_1 , \DDS_0/dds_state_0/N_282 , 
        \DDS_0/dds_state_0/para_9_i_0_1[22] , 
        \DDS_0/dds_state_0/N_459 , \DDS_0/dds_state_0/para_9_i_1[17] , 
        \DDS_0/dds_state_0/N_498 , \DDS_0/dds_state_0/para_9_i_1[21] , 
        \DDS_0/dds_state_0/N_510 , \DDS_0/dds_state_0/para_9_i_1[5] , 
        \DDS_0/dds_state_0/para[5]_net_1 , \DDS_0/dds_state_0/N_319 , 
        \DDS_0/dds_state_0/para_9_i_i_1[7] , 
        \DDS_0/dds_state_0/para[7]_net_1 , \DDS_0/dds_state_0/N_270 , 
        \DDS_0/dds_state_0/N_40 , \DDS_0/dds_state_0/N_269 , 
        \DDS_0/dds_state_0/N_460 , \DDS_0/dds_state_0/N_8 , 
        \DDS_0/dds_state_0/N_273 , \DDS_0/dds_state_0/N_272 , 
        \DDS_0/dds_state_0/N_44 , \DDS_0/dds_state_0/N_277 , 
        \DDS_0/dds_state_0/N_276 , \DDS_0/dds_state_0/N_46 , 
        \DDS_0/dds_state_0/N_281 , \DDS_0/dds_state_0/N_280 , 
        \DDS_0/dds_state_0/N_12 , \DDS_0/dds_state_0/N_285 , 
        \DDS_0/dds_state_0/N_284 , \DDS_0/dds_state_0/N_14 , 
        \DDS_0/dds_state_0/N_289 , \DDS_0/dds_state_0/N_288 , 
        \DDS_0/dds_state_0/N_16 , \DDS_0/dds_state_0/N_293 , 
        \DDS_0/dds_state_0/N_292 , \DDS_0/dds_state_0/N_18 , 
        \DDS_0/dds_state_0/N_297 , \DDS_0/dds_state_0/N_296 , 
        \DDS_0/dds_state_0/N_20 , \DDS_0/dds_state_0/N_301 , 
        \DDS_0/dds_state_0/N_300 , \DDS_0/dds_state_0/N_23 , 
        \DDS_0/dds_state_0/N_305 , \DDS_0/dds_state_0/N_304 , 
        \DDS_0/dds_state_0/N_25 , \DDS_0/dds_state_0/N_310 , 
        \DDS_0/dds_state_0/N_309 , \DDS_0/dds_state_0/N_27 , 
        \DDS_0/dds_state_0/N_314 , \DDS_0/dds_state_0/N_313 , 
        \DDS_0/dds_state_0/N_54 , \DDS_0/dds_state_0/N_318 , 
        \DDS_0/dds_state_0/N_317 , \DDS_0/dds_state_0/N_81 , 
        \DDS_0/dds_state_0/N_323 , \DDS_0/dds_state_0/N_321 , 
        \DDS_0/dds_state_0/N_87 , \DDS_0/dds_state_0/N_328 , 
        \DDS_0/dds_state_0/N_327 , \DDS_0/dds_state_0/N_103 , 
        \DDS_0/dds_state_0/N_333 , \DDS_0/dds_state_0/N_332 , 
        \DDS_0/dds_state_0/N_118 , \DDS_0/dds_state_0/N_337 , 
        \DDS_0/dds_state_0/N_336 , \DDS_0/dds_state_0/N_121 , 
        \DDS_0/dds_state_0/N_464 , \DDS_0/dds_state_0/N_463 , 
        \DDS_0/dds_state_0/N_123 , \DDS_0/dds_state_0/N_468 , 
        \DDS_0/dds_state_0/N_467 , \DDS_0/dds_state_0/N_125 , 
        \DDS_0/dds_state_0/N_472 , \DDS_0/dds_state_0/N_471 , 
        \DDS_0/dds_state_0/N_127 , \DDS_0/dds_state_0/N_476 , 
        \DDS_0/dds_state_0/N_475 , \DDS_0/dds_state_0/N_129 , 
        \DDS_0/dds_state_0/N_480 , \DDS_0/dds_state_0/N_479 , 
        \DDS_0/dds_state_0/N_131 , \DDS_0/dds_state_0/N_484 , 
        \DDS_0/dds_state_0/N_483 , \DDS_0/dds_state_0/N_155 , 
        \DDS_0/dds_state_0/N_488 , \DDS_0/dds_state_0/N_487 , 
        \DDS_0/dds_state_0/N_157 , \DDS_0/dds_state_0/N_492 , 
        \DDS_0/dds_state_0/N_491 , \DDS_0/dds_state_0/N_159 , 
        \DDS_0/dds_state_0/N_496 , \DDS_0/dds_state_0/N_495 , 
        \DDS_0/dds_state_0/N_161 , \DDS_0/dds_state_0/N_500 , 
        \DDS_0/dds_state_0/N_499 , \DDS_0/dds_state_0/N_163 , 
        \DDS_0/dds_state_0/N_504 , \DDS_0/dds_state_0/N_503 , 
        \DDS_0/dds_state_0/N_165 , \DDS_0/dds_state_0/N_508 , 
        \DDS_0/dds_state_0/N_507 , \DDS_0/dds_state_0/N_167 , 
        \DDS_0/dds_state_0/N_512 , \DDS_0/dds_state_0/N_511 , 
        \DDS_0/dds_state_0/N_169 , \DDS_0/dds_state_0/N_516 , 
        \DDS_0/dds_state_0/N_515 , \DDS_0/dds_state_0/N_171 , 
        \DDS_0/dds_state_0/N_518 , \DDS_0/dds_state_0/N_517 , 
        \DDS_0/dds_state_0/N_21 , \DDS_0/dds_state_0/para[0]_net_1 , 
        \DDS_0/dds_state_0/N_223 , \DDS_0/dds_state_0/N_531 , 
        \DDS_0/dds_state_0/N_451 , \DDS_0/dds_state_0/cs[7]_net_1 , 
        \DDS_0/dds_state_0/cs[8]_net_1 , 
        \DDS_0/dds_state_0/fq_ud_RNO_net_1 , 
        \DDS_0/dds_state_0/fq_ud_reg_net_1 , \DDS_0/dds_state_0/N_538 , 
        \DDS_0/dds_state_0/para[22]_net_1 , \DDS_0/dds_state_0/N_535 , 
        \DDS_0/dds_state_0/para_reg[22]_net_1 , 
        \DDS_0/dds_state_0/N_534 , \DDS_0/dds_state_0/para[23]_net_1 , 
        \DDS_0/dds_state_0/para_reg[7]_net_1 , 
        \DDS_0/dds_state_0/para_reg[6]_net_1 , 
        \DDS_0/dds_state_0/para_reg[1]_net_1 , 
        \DDS_0/dds_state_0/para_reg[8]_net_1 , 
        \DDS_0/dds_state_0/para_reg[9]_net_1 , 
        \DDS_0/dds_state_0/para_reg[10]_net_1 , 
        \DDS_0/dds_state_0/para_reg[16]_net_1 , 
        \DDS_0/dds_state_0/para[17]_net_1 , 
        \DDS_0/dds_state_0/para_reg[23]_net_1 , 
        \DDS_0/dds_state_0/para[24]_net_1 , 
        \DDS_0/dds_state_0/para_reg[24]_net_1 , 
        \DDS_0/dds_state_0/para[25]_net_1 , 
        \DDS_0/dds_state_0/para_reg[25]_net_1 , 
        \DDS_0/dds_state_0/para[26]_net_1 , 
        \DDS_0/dds_state_0/para[32]_net_1 , 
        \DDS_0/dds_state_0/para_reg[32]_net_1 , 
        \DDS_0/dds_state_0/para[33]_net_1 , 
        \DDS_0/dds_state_0/para_reg[4]_net_1 , 
        \DDS_0/dds_state_0/para_reg[5]_net_1 , 
        \DDS_0/dds_state_0/para_reg[11]_net_1 , 
        \DDS_0/dds_state_0/para_reg[12]_net_1 , 
        \DDS_0/dds_state_0/para_reg[13]_net_1 , 
        \DDS_0/dds_state_0/para_reg[14]_net_1 , 
        \DDS_0/dds_state_0/para[20]_net_1 , 
        \DDS_0/dds_state_0/para_reg[20]_net_1 , 
        \DDS_0/dds_state_0/para[21]_net_1 , 
        \DDS_0/dds_state_0/para_reg[26]_net_1 , 
        \DDS_0/dds_state_0/para[27]_net_1 , 
        \DDS_0/dds_state_0/para_reg[27]_net_1 , 
        \DDS_0/dds_state_0/para[28]_net_1 , 
        \DDS_0/dds_state_0/para_reg[28]_net_1 , 
        \DDS_0/dds_state_0/para[29]_net_1 , 
        \DDS_0/dds_state_0/para_reg[29]_net_1 , 
        \DDS_0/dds_state_0/para[30]_net_1 , 
        \DDS_0/dds_state_0/para_reg[2]_net_1 , 
        \DDS_0/dds_state_0/para_reg[3]_net_1 , 
        \DDS_0/dds_state_0/para_reg[15]_net_1 , 
        \DDS_0/dds_state_0/para_reg[17]_net_1 , 
        \DDS_0/dds_state_0/para[18]_net_1 , 
        \DDS_0/dds_state_0/para_reg[18]_net_1 , 
        \DDS_0/dds_state_0/para[19]_net_1 , 
        \DDS_0/dds_state_0/para_reg[19]_net_1 , 
        \DDS_0/dds_state_0/para_reg[21]_net_1 , 
        \DDS_0/dds_state_0/para_reg[30]_net_1 , 
        \DDS_0/dds_state_0/para[31]_net_1 , \DDS_0/dds_state_0/N_522 , 
        \DDS_0/dds_state_0/para[34]_net_1 , \DDS_0/dds_state_0/N_524 , 
        \DDS_0/dds_state_0/para[35]_net_1 , \DDS_0/dds_state_0/N_526 , 
        \DDS_0/dds_state_0/para[36]_net_1 , 
        \DDS_0/dds_state_0/para_9[36] , \DDS_0/dds_state_0/N_528 , 
        \DDS_0/dds_state_0/N_224 , \DDS_0/dds_state_0/cs[4]_net_1 , 
        \DDS_0/dds_state_0/cs[5]_net_1 , 
        \DDS_0/dds_state_0/para_1_sqmuxa_1 , 
        \DDS_0/dds_state_0/cs_RNO[3]_net_1 , \DDS_0/dds_state_0/N_227 , 
        \DDS_0/dds_state_0/cs_RNO[4]_net_1 , 
        \DDS_0/dds_state_0/cs[3]_net_1 , 
        \DDS_0/dds_state_0/cs_RNO[6]_net_1 , \DDS_0/dds_state_0/N_80 , 
        \DDS_0/dds_state_0/N_226 , \DDS_0/dds_state_0/cs_RNO[8]_net_1 , 
        \DDS_0/dds_state_0/w_clk_RNO_net_1 , 
        \DDS_0/dds_state_0/reset_RNO_net_1 , 
        \DDS_0/dds_state_0/cs[1]_net_1 , 
        \DDS_0/dds_state_0/para_9[33] , \DDS_0/dds_state_0/para_9[34] , 
        \DDS_0/dds_state_0/para_9[35] , \DDS_0/dds_state_0/N_203 , 
        \DDS_0/dds_state_0/N_38 , \DDS_0/dds_state_0/N_228 , 
        \DDS_0/dds_state_0/N_225 , \DDS_0/dds_state_0/cs_RNO[5]_net_1 , 
        \DDS_0/dds_state_0/fq_ud_reg_RNO_net_1 , 
        \DDS_0/dds_state_0/w_clk_reg_RNO_net_1 , 
        \DDS_0/dds_state_0/cs_RNO[1]_net_1 , 
        \DDS_0/dds_state_0/cs_i[0]_net_1 , \DDS_0/dds_state_0/N_229 , 
        \DDS_0/dds_state_0/state_over_RNO_net_1 , 
        \DDS_0/dds_state_0/cs[6]_net_1 , 
        \DDS_0/dds_state_0/cs[2]_net_1 , 
        \DDS_0/dds_coder_0/m12_2_net_1 , 
        \DDS_0/dds_coder_0/m12_0_net_1 , \DDS_0/dds_coder_0/m8_2 , 
        \DDS_0/dds_coder_0/m8_1 , \DDS_0/dds_coder_0/m3_e_1_net_1 , 
        \DDS_0/dds_coder_0/i_RNO[3]_net_1 , 
        \DDS_0/dds_coder_0/N_18_mux , 
        \DDS_0/dds_coder_0/i_RNO[0]_net_1 , 
        \DDS_0/dds_coder_0/i_RNO[2]_net_1 , 
        \DDS_0/dds_coder_0/i_RNO[1]_net_1 , \timer_top_0/dataout[0] , 
        \timer_top_0/dataout[1] , \timer_top_0/dataout[2] , 
        \timer_top_0/dataout[3] , \timer_top_0/dataout[4] , 
        \timer_top_0/dataout[5] , \timer_top_0/dataout[6] , 
        \timer_top_0/dataout[7] , \timer_top_0/dataout[8] , 
        \timer_top_0/dataout[9] , \timer_top_0/dataout[10] , 
        \timer_top_0/dataout[11] , \timer_top_0/dataout[12] , 
        \timer_top_0/dataout[13] , \timer_top_0/dataout[14] , 
        \timer_top_0/dataout[15] , \timer_top_0/dataout[16] , 
        \timer_top_0/dataout[17] , \timer_top_0/dataout[18] , 
        \timer_top_0/dataout[19] , \timer_top_0/dataout[20] , 
        \timer_top_0/dataout[21] , \timer_top_0/timer_0_time_up , 
        \timer_top_0/state_switch_0_state_start , 
        \timer_top_0/state_switch_0_state_over_n , 
        \timer_top_0/timer_0/timedata[1]_net_1 , 
        \timer_top_0/timer_0/timedata[0]_net_1 , 
        \timer_top_0/timer_0/timedata[3]_net_1 , 
        \timer_top_0/timer_0/DWACT_FINC_E[0] , 
        \timer_top_0/timer_0/timedata[8]_net_1 , 
        \timer_top_0/timer_0/DWACT_FINC_E[4] , 
        \timer_top_0/timer_0/DWACT_FINC_E[7] , 
        \timer_top_0/timer_0/DWACT_FINC_E[6] , 
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 , 
        \timer_top_0/timer_0/timedata_4[1] , 
        \timer_top_0/timer_0/I_5_2 , 
        \timer_top_0/timer_0/timedata_4[2] , 
        \timer_top_0/timer_0/I_7_2 , 
        \timer_top_0/timer_0/timedata_4[3] , 
        \timer_top_0/timer_0/I_9_2 , 
        \timer_top_0/timer_0/timedata_4[4] , 
        \timer_top_0/timer_0/I_12_2 , 
        \timer_top_0/timer_0/timedata_4[5] , 
        \timer_top_0/timer_0/I_14_1 , 
        \timer_top_0/timer_0/timedata_4[6] , 
        \timer_top_0/timer_0/I_17_0 , 
        \timer_top_0/timer_0/timedata_4[7] , 
        \timer_top_0/timer_0/I_20_0 , 
        \timer_top_0/timer_0/timedata_4[8] , 
        \timer_top_0/timer_0/I_23_0 , 
        \timer_top_0/timer_0/timedata_4[9] , 
        \timer_top_0/timer_0/I_26_0 , 
        \timer_top_0/timer_0/timedata_4[10] , 
        \timer_top_0/timer_0/I_28_0 , 
        \timer_top_0/timer_0/timedata_4[11] , 
        \timer_top_0/timer_0/I_32_2 , 
        \timer_top_0/timer_0/timedata_4[12] , 
        \timer_top_0/timer_0/I_35_1 , 
        \timer_top_0/timer_0/timedata_4[13] , 
        \timer_top_0/timer_0/I_37_1 , 
        \timer_top_0/timer_0/timedata_4[14] , 
        \timer_top_0/timer_0/I_40 , 
        \timer_top_0/timer_0/timedata_4[15] , 
        \timer_top_0/timer_0/I_43 , 
        \timer_top_0/timer_0/timedata_4[16] , 
        \timer_top_0/timer_0/I_46 , 
        \timer_top_0/timer_0/timedata_4[17] , 
        \timer_top_0/timer_0/I_49 , 
        \timer_top_0/timer_0/timedata_4[18] , 
        \timer_top_0/timer_0/I_53 , 
        \timer_top_0/timer_0/timedata_4[19] , 
        \timer_top_0/timer_0/I_56 , 
        \timer_top_0/timer_0/timedata_4[20] , 
        \timer_top_0/timer_0/I_59 , 
        \timer_top_0/timer_0/timedata_4[21] , 
        \timer_top_0/timer_0/I_62 , 
        \timer_top_0/timer_0/timedata_4[0] , 
        \timer_top_0/timer_0/time_up_RNO_net_1 , 
        \timer_top_0/timer_0/cmp_result , 
        \timer_top_0/timer_0/timedata[2]_net_1 , 
        \timer_top_0/timer_0/timedata[4]_net_1 , 
        \timer_top_0/timer_0/timedata[5]_net_1 , 
        \timer_top_0/timer_0/timedata[6]_net_1 , 
        \timer_top_0/timer_0/timedata[7]_net_1 , 
        \timer_top_0/timer_0/timedata[9]_net_1 , 
        \timer_top_0/timer_0/timedata[10]_net_1 , 
        \timer_top_0/timer_0/timedata[11]_net_1 , 
        \timer_top_0/timer_0/timedata[12]_net_1 , 
        \timer_top_0/timer_0/timedata[13]_net_1 , 
        \timer_top_0/timer_0/timedata[14]_net_1 , 
        \timer_top_0/timer_0/timedata[15]_net_1 , 
        \timer_top_0/timer_0/timedata[16]_net_1 , 
        \timer_top_0/timer_0/timedata[17]_net_1 , 
        \timer_top_0/timer_0/timedata[18]_net_1 , 
        \timer_top_0/timer_0/timedata[19]_net_1 , 
        \timer_top_0/timer_0/timedata[20]_net_1 , 
        \timer_top_0/timer_0/timedata[21]_net_1 , 
        \timer_top_0/timer_0/N_2 , 
        \timer_top_0/timer_0/DWACT_FINC_E[28] , 
        \timer_top_0/timer_0/DWACT_FINC_E[13] , 
        \timer_top_0/timer_0/DWACT_FINC_E[15] , 
        \timer_top_0/timer_0/N_3 , 
        \timer_top_0/timer_0/DWACT_FINC_E[14] , 
        \timer_top_0/timer_0/N_4 , 
        \timer_top_0/timer_0/DWACT_FINC_E[9] , 
        \timer_top_0/timer_0/DWACT_FINC_E[12] , 
        \timer_top_0/timer_0/N_5 , 
        \timer_top_0/timer_0/DWACT_FINC_E[10] , 
        \timer_top_0/timer_0/DWACT_FINC_E[2] , 
        \timer_top_0/timer_0/DWACT_FINC_E[5] , 
        \timer_top_0/timer_0/N_6 , 
        \timer_top_0/timer_0/DWACT_FINC_E[11] , 
        \timer_top_0/timer_0/N_7 , \timer_top_0/timer_0/N_8 , 
        \timer_top_0/timer_0/N_9 , 
        \timer_top_0/timer_0/DWACT_FINC_E[8] , 
        \timer_top_0/timer_0/N_10 , \timer_top_0/timer_0/N_12 , 
        \timer_top_0/timer_0/N_13 , 
        \timer_top_0/timer_0/DWACT_FINC_E[3] , 
        \timer_top_0/timer_0/N_15 , \timer_top_0/timer_0/N_16 , 
        \timer_top_0/timer_0/N_17 , 
        \timer_top_0/timer_0/DWACT_FINC_E[1] , 
        \timer_top_0/timer_0/N_18 , \timer_top_0/timer_0/N_20 , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_10_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_7_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_7_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_19_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_23_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_21_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_6_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_7_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_6_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_7_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_11_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_8_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_11_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_8_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_7_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_27_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_6_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_24_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_20_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR2A_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_17_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_26_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_13_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_9_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_14_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_10_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_12_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_10_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_6_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_8_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_16_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_8_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_10_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_28_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_4_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_8_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_22_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_9_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_5_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_9_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_18_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_9_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_12_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_6_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_11_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AO1D_0_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_9_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_2_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_3_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_1_Y , 
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_1_Y , 
        \timer_top_0/state_switch_0/clk_en_scale_0_0_a6_0_a5_net_1 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[10] , 
        \timer_top_0/state_switch_0/N_252 , 
        \timer_top_0/state_switch_0/N_254 , 
        \timer_top_0/state_switch_0/N_253 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[14] , 
        \timer_top_0/state_switch_0/N_262 , 
        \timer_top_0/state_switch_0/N_264 , 
        \timer_top_0/state_switch_0/N_263 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[9] , 
        \timer_top_0/state_switch_0/N_202 , 
        \timer_top_0/state_switch_0/N_204 , 
        \timer_top_0/state_switch_0/N_203 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[8] , 
        \timer_top_0/state_switch_0/N_247 , 
        \timer_top_0/state_switch_0/N_249 , 
        \timer_top_0/state_switch_0/N_248 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[0] , 
        \timer_top_0/state_switch_0/N_242 , 
        \timer_top_0/state_switch_0/N_244 , 
        \timer_top_0/state_switch_0/N_243 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[15] , 
        \timer_top_0/state_switch_0/N_187 , 
        \timer_top_0/state_switch_0/N_189 , 
        \timer_top_0/state_switch_0/N_188 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[12] , 
        \timer_top_0/state_switch_0/N_257 , 
        \timer_top_0/state_switch_0/N_259 , 
        \timer_top_0/state_switch_0/N_258 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[13] , 
        \timer_top_0/state_switch_0/N_192 , 
        \timer_top_0/state_switch_0/N_194 , 
        \timer_top_0/state_switch_0/N_193 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[4] , 
        \timer_top_0/state_switch_0/N_222 , 
        \timer_top_0/state_switch_0/N_224 , 
        \timer_top_0/state_switch_0/N_223 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[11] , 
        \timer_top_0/state_switch_0/N_197 , 
        \timer_top_0/state_switch_0/N_199 , 
        \timer_top_0/state_switch_0/N_198 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[1] , 
        \timer_top_0/state_switch_0/N_237 , 
        \timer_top_0/state_switch_0/N_239 , 
        \timer_top_0/state_switch_0/N_238 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[5] , 
        \timer_top_0/state_switch_0/N_217 , 
        \timer_top_0/state_switch_0/N_219 , 
        \timer_top_0/state_switch_0/N_218 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[6] , 
        \timer_top_0/state_switch_0/N_212 , 
        \timer_top_0/state_switch_0/N_214 , 
        \timer_top_0/state_switch_0/N_213 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[7] , 
        \timer_top_0/state_switch_0/N_207 , 
        \timer_top_0/state_switch_0/N_209 , 
        \timer_top_0/state_switch_0/N_208 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[2] , 
        \timer_top_0/state_switch_0/N_232 , 
        \timer_top_0/state_switch_0/N_234 , 
        \timer_top_0/state_switch_0/N_233 , 
        \timer_top_0/state_switch_0/dataout_0_0_0_1[3] , 
        \timer_top_0/state_switch_0/N_227 , 
        \timer_top_0/state_switch_0/N_229 , 
        \timer_top_0/state_switch_0/N_228 , 
        \timer_top_0/state_switch_0/state_over_n_0_i_0 , 
        \timer_top_0/state_switch_0/N_297 , 
        \timer_top_0/state_switch_0/N_280 , 
        \timer_top_0/state_switch_0/state_start5_0_0_1 , 
        \timer_top_0/state_switch_0/N_289 , 
        \timer_top_0/state_switch_0/N_168 , 
        \timer_top_0/state_switch_0/state_start5_0_0_a2_1_0_net_1 , 
        \timer_top_0/state_switch_0/state_start5_0_0_a2_2_0_net_1 , 
        \timer_top_0/state_switch_0/state_start5_0_0_a2_0_0 , 
        \timer_top_0/state_switch_0/N_295 , 
        \timer_top_0/state_switch_0/N_284 , 
        \timer_top_0/state_switch_0/dataout_RNO[3]_net_1 , 
        \timer_top_0/state_switch_0/N_225 , 
        \timer_top_0/state_switch_0/N_226 , 
        \timer_top_0/state_switch_0/N_285 , 
        \timer_top_0/state_switch_0/N_293 , 
        \timer_top_0/state_switch_0/dataout_RNO[9]_net_1 , 
        \timer_top_0/state_switch_0/N_200 , 
        \timer_top_0/state_switch_0/N_201 , 
        \timer_top_0/state_switch_0/N_282 , 
        \timer_top_0/state_switch_0/N_78 , 
        \timer_top_0/state_switch_0/N_278 , 
        \timer_top_0/state_switch_0/N_279 , 
        \timer_top_0/state_switch_0/dataout_RNO[11]_net_1 , 
        \timer_top_0/state_switch_0/N_195 , 
        \timer_top_0/state_switch_0/N_196 , 
        \timer_top_0/state_switch_0/state_start5 , 
        \timer_top_0/state_switch_0/N_296 , 
        \timer_top_0/state_switch_0/dataout_RNO[13]_net_1 , 
        \timer_top_0/state_switch_0/N_190 , 
        \timer_top_0/state_switch_0/N_191 , 
        \timer_top_0/state_switch_0/dataout_RNO[15]_net_1 , 
        \timer_top_0/state_switch_0/N_185 , 
        \timer_top_0/state_switch_0/N_186 , 
        \timer_top_0/state_switch_0/dataout_RNO[7]_net_1 , 
        \timer_top_0/state_switch_0/N_205 , 
        \timer_top_0/state_switch_0/N_206 , 
        \timer_top_0/state_switch_0/dataout_RNO[6]_net_1 , 
        \timer_top_0/state_switch_0/N_210 , 
        \timer_top_0/state_switch_0/N_211 , 
        \timer_top_0/state_switch_0/dataout_RNO[5]_net_1 , 
        \timer_top_0/state_switch_0/N_215 , 
        \timer_top_0/state_switch_0/N_216 , 
        \timer_top_0/state_switch_0/dataout_RNO[4]_net_1 , 
        \timer_top_0/state_switch_0/N_220 , 
        \timer_top_0/state_switch_0/N_221 , 
        \timer_top_0/state_switch_0/dataout_RNO[2]_net_1 , 
        \timer_top_0/state_switch_0/N_230 , 
        \timer_top_0/state_switch_0/N_231 , 
        \timer_top_0/state_switch_0/dataout_RNO[1]_net_1 , 
        \timer_top_0/state_switch_0/N_235 , 
        \timer_top_0/state_switch_0/N_236 , 
        \timer_top_0/state_switch_0/dataout_RNO[0]_net_1 , 
        \timer_top_0/state_switch_0/N_240 , 
        \timer_top_0/state_switch_0/N_241 , 
        \timer_top_0/state_switch_0/dataout_RNO[8]_net_1 , 
        \timer_top_0/state_switch_0/N_245 , 
        \timer_top_0/state_switch_0/N_246 , 
        \timer_top_0/state_switch_0/dataout_RNO[10]_net_1 , 
        \timer_top_0/state_switch_0/N_250 , 
        \timer_top_0/state_switch_0/N_251 , 
        \timer_top_0/state_switch_0/dataout_RNO[12]_net_1 , 
        \timer_top_0/state_switch_0/N_255 , 
        \timer_top_0/state_switch_0/N_256 , 
        \timer_top_0/state_switch_0/dataout_RNO[14]_net_1 , 
        \timer_top_0/state_switch_0/N_260 , 
        \timer_top_0/state_switch_0/N_261 , 
        \timer_top_0/state_switch_0/dataout_RNO[21]_net_1 , 
        \timer_top_0/state_switch_0/dataout_RNO[20]_net_1 , 
        \timer_top_0/state_switch_0/N_266 , 
        \timer_top_0/state_switch_0/N_268 , 
        \timer_top_0/state_switch_0/N_270 , 
        \timer_top_0/state_switch_0/clk_en_st1ms_RNO_net_1 , 
        \timer_top_0/state_switch_0/clk_en_scan_RNO_net_1 , 
        \timer_top_0/state_switch_0/clk_en_noise_RNO_net_1 , 
        \timer_top_0/state_switch_0/dataout_RNO[16]_net_1 , 
        \timer_top_0/state_switch_0/dataout_RNO[17]_net_1 , 
        \timer_top_0/state_switch_0/dataout_RNO[18]_net_1 , 
        \timer_top_0/state_switch_0/clk_en_pluse_RNO_net_1 , 
        \timer_top_0/state_switch_0/dataout_RNO[19]_net_1 , 
        \timer_top_0/state_switch_0/N_272 , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[1] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[2] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[3] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[4] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[5] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[6] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[7] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[8] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[9] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[10] , 
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[11] , 
        \Signal_Noise_Acq_0/signal_data_t[4] , 
        \Signal_Noise_Acq_0/signal_data_t[5] , 
        \Signal_Noise_Acq_0/signal_data_t[6] , 
        \Signal_Noise_Acq_0/signal_data_t[7] , 
        \Signal_Noise_Acq_0/signal_data_t[8] , 
        \Signal_Noise_Acq_0/signal_data_t[9] , 
        \Signal_Noise_Acq_0/signal_data_t[10] , 
        \Signal_Noise_Acq_0/signal_data_t[11] , 
        \Signal_Noise_Acq_0/signal_data_t[12] , 
        \Signal_Noise_Acq_0/signal_data_t[13] , 
        \Signal_Noise_Acq_0/signal_data_t[14] , 
        \Signal_Noise_Acq_0/signal_data_t[15] , 
        \Signal_Noise_Acq_0/un1_signal_acq_0[0] , 
        \Signal_Noise_Acq_0/un1_signal_acq_0[1] , 
        \Signal_Noise_Acq_0/un1_signal_acq_0[2] , 
        \Signal_Noise_Acq_0/un1_signal_acq_0[3] , 
        \Signal_Noise_Acq_0/signal_acq_0_Signal_acq_clk , 
        \Signal_Noise_Acq_0/MX2_RD_0_inst , 
        \Signal_Noise_Acq_0/MX2_RD_2_inst , 
        \Signal_Noise_Acq_0/n_adc_1_10 , 
        \Signal_Noise_Acq_0/n_adc_1_9 , \Signal_Noise_Acq_0/n_adc_1_8 , 
        \Signal_Noise_Acq_0/n_adc_1_7 , \Signal_Noise_Acq_0/n_adc_1_6 , 
        \Signal_Noise_Acq_0/n_adc_1_5 , \Signal_Noise_Acq_0/n_adc_1_4 , 
        \Signal_Noise_Acq_0/n_adc_1_3 , \Signal_Noise_Acq_0/n_adc_1_2 , 
        \Signal_Noise_Acq_0/n_adc_1_1 , \Signal_Noise_Acq_0/n_adc_1_0 , 
        \Signal_Noise_Acq_0/n_adc_1 , 
        \Signal_Noise_Acq_0/MX2_RD_4_inst , 
        \Signal_Noise_Acq_0/MX2_RD_5_inst , 
        \Signal_Noise_Acq_0/MX2_RD_7_inst , 
        \Signal_Noise_Acq_0/MX2_RD_6_inst , 
        \Signal_Noise_Acq_0/MX2_RD_11_inst , 
        \Signal_Noise_Acq_0/MX2_RD_1_inst , 
        \Signal_Noise_Acq_0/MX2_RD_9_inst , 
        \Signal_Noise_Acq_0/MX2_RD_3_inst , 
        \Signal_Noise_Acq_0/MX2_RD_10_inst , 
        \Signal_Noise_Acq_0/MX2_RD_8_inst , 
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout , 
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add , 
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree , 
        \Signal_Noise_Acq_0/signal_acq_0/clkout , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[13] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[14] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[15] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[17] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[18] , 
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[19] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone , 
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/addrout[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/addrout[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/addrout[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[9] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[11] , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_1_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/ADD_20x20_slow_I19_Y_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_38_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_40_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m41_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m42_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m43_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m44_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m45_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m46_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m47_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m70_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_RNO_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_1_sqmuxa , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_313 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_311 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_6_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_7_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_8_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_9_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_10_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_11_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_12_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_13_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_14_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_15_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_16_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_17_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_18_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_19_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_20 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_21 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_22 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_23 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_24 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_25 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_26 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_27 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_28 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_29 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_30 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_31 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_32 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_33 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_34 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_35 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_37 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_38 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_39 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_40 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_41 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_42 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_43 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_44 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_45 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_46 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_47 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_48 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_49 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_50 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_51 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_52 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_53 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_54 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_55 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_56 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_57 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_58 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_59 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_60 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_61 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_62 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_63 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_64 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_65 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_66 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_69 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_70 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_71 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_72 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_73 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_74 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_75 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_76 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_77 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_78 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_79 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_80 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_81 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_82 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_84 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_85 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_86 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_87 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_88 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_89 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_90 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_91 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_92 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_93 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_94 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_95 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_96 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_97 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_99 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_100 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_101 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_102 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_103 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_104 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_105 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_106 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_107 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_108 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_109 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_110 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_111 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_112 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_114 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_115 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_116 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_117 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_118 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_119 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_120 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_121 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_122 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_123 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_124 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_125 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_126 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_127 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_128 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_129 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_130 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_131 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_132 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_133 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_134 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_135 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_136 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_137 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_138 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_139 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_140 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_141 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_142 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_143 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_145 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_146 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_147 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_148 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_149 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_150 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_151 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_152 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_153 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_154 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_155 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_156 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_157 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_158 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_159 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_160 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_161 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_162 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_163 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_164 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_165 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_166 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_167 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_168 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_169 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_170 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_171 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_172 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_173 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_174 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_176 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_177 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_178 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_179 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_180 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_181 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_182 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_183 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_184 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_185 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_186 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_187 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_188 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_189 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_191 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_192 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_193 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_194 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_195 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_196 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_197 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_198 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_199 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_200 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_201 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_202 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_203 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_204 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_206 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_207 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_208 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_209 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_210 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_211 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_212 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_213 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_214 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_215 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_216 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_217 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_218 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_219 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_221 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_222 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_223 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_224 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_225 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_226 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_227 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_228 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_229 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_230 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_231 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_232 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_233 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_234 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_236 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_237 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_238 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_239 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_240 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_241 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_242 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_243 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_244 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_245 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_246 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_247 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_248 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_249 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_251 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_252 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_253 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_254 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_255 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_256 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_257 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_258 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_259 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_260 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_261 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_262 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_263 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_264 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_266 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_267 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_268 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_269 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_270 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_271 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_272 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_273 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_274 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_275 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_276 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_277 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_278 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_279 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_281 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_282 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_283 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_284 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_285 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_286 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_287 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_288 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_289 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_290 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_291 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_292 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_293 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_294 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_296 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_297 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_298 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_299 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_300 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_301 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_302 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_303 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_304 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_305 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_306 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_307 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_308 , 
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_309 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/clk_add_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_12 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_0_i_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_8_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_9 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_8_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_7 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_11 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_12 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_10_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_9_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_11 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_7 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_10 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_10 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_9 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_20 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_11 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_12_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_26 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_5 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_1_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[1]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N142 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[3]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N168 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N160 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_65 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I0_un1_CO1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[2]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I2_un1_CO1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N146 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I4_un1_CO1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N152 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I6_un1_CO1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I10_un1_CO1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[1]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[2]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[3]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[4]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[5]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[6]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[7]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_48_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[8]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_46_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[9]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_44_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[10]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_42_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[11]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/entop_RNO_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[14]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[15]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[13]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m38 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m39 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c2 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c4 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c10 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c12 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c14 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNO_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_RNO_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n2 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n3 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n4 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n5 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n7 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n9 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n10 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n11 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n12 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n13 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n14 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n15 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_10_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_5_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[10] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[7] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[8] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[6] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[4] , 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[5] , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/ADD_20x20_slow_I19_Y_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m41_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m42_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m43_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m44_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m45_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m46_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m47_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m70_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/ADD_20x20_slow_I19_Y_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m41_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m42_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m43_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m44_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m45_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m46_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m47_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m70_6 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/ADD_20x20_slow_I19_Y_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m41_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m42_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m43_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m44_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m45_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m46_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m47_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m70_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/ADD_20x20_slow_I19_Y_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_38_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m41_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m42_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m43_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m44_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m45_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m46_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m47_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m70_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/ADD_20x20_slow_I19_Y_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_38_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m41_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m42_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m43_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m44_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m45_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m46_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m47_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m70_3 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[1]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[3]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIKJJB2[2]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNILKJB2[3]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[0]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[2]_net_1 , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[0] , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[1] , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[2] , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[3] , 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/N_2 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/ADD_20x20_slow_I19_Y , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m41 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m42 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m43 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m44 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m45 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m46 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m47 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m70 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_70_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_2_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_68_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i2_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_66_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i4_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_64_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i6_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_62_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i8_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_60_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i10_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_58_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i12_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_56_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i14_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_54_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i16_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_52_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i18_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_50_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i20_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/ADD_20x20_slow_I19_Y_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_41_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_37_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i22_mux , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_39_i , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m41_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m42_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m43_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m44_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m45_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m46_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m47_4 , 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m70_4 , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[7] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0_en , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[6] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[7] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] , 
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk_RNO_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/un1_clk_wire , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_RNO_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_RNO_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/un1_noise_addr_0_i[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n7 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n5 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n11 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/DWACT_FINC_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[2]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i6_mux , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_1_sqmuxa , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_11 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_14_i , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_i , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_12_i , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i2_mux , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10_i , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i4_mux , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_5_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_7_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_9_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_12_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_41 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[0]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[1]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[3]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[4]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[0]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[1]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[2]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[3]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[4]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_11 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_7 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_5 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3_0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_4_0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/en_RNO_0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_e0 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n11 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n5 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n7 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[0]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[1]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[2]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[3]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[4]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[7]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]_net_1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[6] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[10] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[7] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[8] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[5] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[3] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[5] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_11 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_7 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_5 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[4] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_149_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_75_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_127_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_140_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_14_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_147_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_144_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_13_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_1_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_162_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_22_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_111_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_126_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_85_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_16_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_3_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_167_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_165_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_34_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_122_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_118_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_94_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_129_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_17_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_13_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_137_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_11_net , GND, 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_7_net , VCC, 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_18_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_138_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_19_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_99_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_161_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_108_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_47_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_73_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_21_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_101_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_81_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_135_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_28_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_89_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_87_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_74_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_39_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_53_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_8_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_12_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_64_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_103_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_59_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_120_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_145_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_4_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_104_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_50_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_97_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_43_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_79_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_151_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_69_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_106_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_46_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_78_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_31_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_153_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_55_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_128_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_48_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_113_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_136_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_24_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_139_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_84_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_130_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_142_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_70_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_134_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_156_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_102_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_71_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_37_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_29_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_51_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_83_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_33_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_42_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_160_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_15_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_15_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_164_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_10_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_77_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_163_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_157_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_93_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_9_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_119_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_57_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_116_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_98_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_27_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_13_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_152_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_65_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_67_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_96_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_15_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_107_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_112_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_7_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_132_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_82_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_36_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_124_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_63_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_150_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_95_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_6_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_146_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_100_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_76_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_60_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_38_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_121_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_11_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_41_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_45_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_56_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_66_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_131_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_72_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_148_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_158_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_80_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_166_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_92_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_125_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_40_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_20_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_52_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_14_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_14_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_32_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_105_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_68_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_117_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_23_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_10_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_2_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_61_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_62_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_26_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_109_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_133_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_141_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_143_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_0_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_159_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_54_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_90_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_154_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_30_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_91_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_8_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_110_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_5_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_114_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_123_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_35_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_49_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_86_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_6_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_12_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_25_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_155_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_88_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_58_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_7_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_115_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_3_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_4_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_2_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_5_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_9_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_12_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_44_Y , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_11_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_0_net , 
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_1_net , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/un1_noise_addr_1_i[0] , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n9 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n8 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n7 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n6 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n5 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n4 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n3 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n2 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n1 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c10 , 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n11 , 
        \bri_dump_sw_0/reset_out_0_net_1 , 
        \bri_dump_sw_0/dump_start_5 , 
        \bri_dump_sw_0/reset_out_5_net_1 , 
        \bri_dump_sw_0/dump_start_RNO_net_1 , 
        \bri_dump_sw_0/pluse_start_5 , 
        \bri_dump_sw_0/pluse_start_RNO_net_1 , 
        \bri_dump_sw_0/off_test_5 , \bri_dump_sw_0/phase_ctr_5 , 
        \bri_dump_sw_0/phase_ctr_RNO_net_1 , 
        \bri_dump_sw_0/off_test_RNO_net_1 , 
        \bri_dump_sw_0/turn_delay_4 , 
        \bri_dump_sw_0/dumpoff_ctr_RNO_net_1 , 
        \bri_dump_sw_0/dumpoff_ctr_5 , 
        \bri_dump_sw_0/tetw_pluse_RNO_net_1 , 
        \bri_dump_sw_0/tetw_pluse_5 , \CAL_0/cal_para_out[0] , 
        \CAL_0/cal_para_out[1] , \CAL_0/cal_para_out[2] , 
        \CAL_0/cal_para_out[3] , \CAL_0/cal_para_out[4] , 
        \CAL_0/cal_para_out[5] , \CAL_0/cal_div_0/count[1]_net_1 , 
        \CAL_0/cal_div_0/count[0]_net_1 , 
        \CAL_0/cal_div_0/count[3]_net_1 , 
        \CAL_0/cal_div_0/DWACT_FINC_E[0] , 
        \CAL_0/cal_div_0/clear_n4_NE_2 , \CAL_0/cal_div_0/clear_n4_0 , 
        \CAL_0/cal_div_0/clear_n4_NE_1 , 
        \CAL_0/cal_div_0/count[2]_net_1 , \CAL_0/cal_div_0/clear_n4_3 , 
        \CAL_0/cal_div_0/clear_n4_NE_0 , 
        \CAL_0/cal_div_0/count[5]_net_1 , \CAL_0/cal_div_0/clear_n4_4 , 
        \CAL_0/cal_div_0/clear_n , \CAL_0/cal_div_0/count_5[1] , 
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 , \CAL_0/cal_div_0/I_5 , 
        \CAL_0/cal_div_0/count_5[2] , \CAL_0/cal_div_0/I_7 , 
        \CAL_0/cal_div_0/count_5[3] , \CAL_0/cal_div_0/I_9 , 
        \CAL_0/cal_div_0/count_5[4] , \CAL_0/cal_div_0/I_12 , 
        \CAL_0/cal_div_0/count_5[5] , \CAL_0/cal_div_0/I_14 , 
        \CAL_0/cal_div_0/count_5[0] , \CAL_0/cal_div_0/N_35 , 
        \CAL_0/cal_div_0/cal_RNO_net_1 , 
        \CAL_0/cal_div_0/count[4]_net_1 , \CAL_0/cal_div_0/N_2 , 
        \CAL_0/cal_div_0/N_4 , \PLUSE_0/i_9[0] , \PLUSE_0/i_9[1] , 
        \PLUSE_0/i_4[2] , \PLUSE_0/i_4[3] , 
        \PLUSE_0/qq_state_0_stateover , \PLUSE_0/qq_para3[0] , 
        \PLUSE_0/qq_para3[1] , \PLUSE_0/qq_para3[2] , 
        \PLUSE_0/qq_para3[3] , \PLUSE_0/qq_para3[4] , 
        \PLUSE_0/qq_para3[5] , \PLUSE_0/qq_para2[0] , 
        \PLUSE_0/qq_para2[1] , \PLUSE_0/qq_para2[2] , 
        \PLUSE_0/qq_para2[3] , \PLUSE_0/qq_para2[4] , 
        \PLUSE_0/qq_para2[5] , \PLUSE_0/qq_para1[0] , 
        \PLUSE_0/qq_para1[1] , \PLUSE_0/qq_para1[2] , 
        \PLUSE_0/qq_para1[3] , \PLUSE_0/count_9[0] , 
        \PLUSE_0/count_9[1] , \PLUSE_0/count_9[2] , 
        \PLUSE_0/count_9[3] , \PLUSE_0/count_9[4] , \PLUSE_0/up , 
        \PLUSE_0/count_8[0] , \PLUSE_0/count_8[1] , 
        \PLUSE_0/count_8[2] , \PLUSE_0/count_8[3] , 
        \PLUSE_0/count_8[4] , \PLUSE_0/count_2[5] , 
        \PLUSE_0/count_2[6] , \PLUSE_0/count_2[7] , 
        \PLUSE_0/bri_coder_0_half , \PLUSE_0/half_para[0] , 
        \PLUSE_0/half_para[1] , \PLUSE_0/half_para[2] , 
        \PLUSE_0/half_para[3] , \PLUSE_0/half_para[4] , 
        \PLUSE_0/half_para[5] , \PLUSE_0/half_para[6] , 
        \PLUSE_0/half_para[7] , \PLUSE_0/i_1[4] , \PLUSE_0/i_3[2] , 
        \PLUSE_0/i_3[3] , \PLUSE_0/i_8[0] , \PLUSE_0/i_8[1] , 
        \PLUSE_0/i_7[0] , \PLUSE_0/i_7[1] , \PLUSE_0/i_2[2] , 
        \PLUSE_0/i_2[3] , \PLUSE_0/qq_state_1_stateover , 
        \PLUSE_0/count_7[0] , \PLUSE_0/count_7[1] , 
        \PLUSE_0/count_7[2] , \PLUSE_0/count_7[3] , 
        \PLUSE_0/count_7[4] , \PLUSE_0/down , 
        \PLUSE_0/qq_state_0/cs_RNO_1[2]_net_1 , 
        \PLUSE_0/qq_state_0/cs4 , \PLUSE_0/qq_state_0/N_89 , 
        \PLUSE_0/qq_state_0/N_88 , 
        \PLUSE_0/qq_state_0/cs_RNO_1[3]_net_1 , 
        \PLUSE_0/qq_state_0/N_86 , \PLUSE_0/qq_state_0/N_87 , 
        \PLUSE_0/qq_state_0/Q1Q8_Q2Q7_RNO_net_1 , 
        \PLUSE_0/qq_state_0/N_79 , \PLUSE_0/qq_state_0/cs[4]_net_1 , 
        \PLUSE_0/qq_state_0/stateover_RNO_0 , 
        \PLUSE_0/qq_state_0/N_84 , \PLUSE_0/qq_state_0/N_82 , 
        \PLUSE_0/qq_state_0/cs[1]_net_1 , 
        \PLUSE_0/qq_state_0/cs[3]_net_1 , 
        \PLUSE_0/qq_state_0/cs_RNO_2[4] , 
        \PLUSE_0/qq_state_0/cs_RNO_1[1] , 
        \PLUSE_0/qq_state_0/cs_i[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_0_4[1] , \PLUSE_0/qq_coder_0/i_0_1[1] , 
        \PLUSE_0/qq_coder_0/i_0_2[1] , \PLUSE_0/qq_coder_0/i_0_0[1] , 
        \PLUSE_0/qq_coder_0/un1_count_1[0] , 
        \PLUSE_0/qq_coder_0/i_reg10_NE_3[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_2[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_3[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_NE_0[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_NE_2[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_0[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_2[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_0[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_1[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_2[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_0[0]_net_1 , 
        \PLUSE_0/qq_coder_0/i_reg10_NE[0]_net_1 , 
        \PLUSE_0/qq_coder_0/un1_qq_para2_i[0] , 
        \PLUSE_0/qq_coder_0/i_RNO_2[2] , 
        \PLUSE_0/qq_coder_0/i_RNO_6[1] , 
        \PLUSE_0/qq_coder_0/i_RNO_7[0] , 
        \PLUSE_0/qq_coder_0/i_RNO_2[3] , 
        \PLUSE_0/bri_timer_0/clken_net_1 , 
        \PLUSE_0/bri_timer_0/count_e0 , \PLUSE_0/bri_timer_0/count_n7 , 
        \PLUSE_0/bri_timer_0/count_c5 , \PLUSE_0/bri_timer_0/count_c4 , 
        \PLUSE_0/bri_timer_0/count_n1 , \PLUSE_0/bri_timer_0/count_n5 , 
        \PLUSE_0/bri_timer_0/count_n6 , \PLUSE_0/bri_timer_0/count_n4 , 
        \PLUSE_0/bri_timer_0/count_c2 , \PLUSE_0/bri_timer_0/count_n3 , 
        \PLUSE_0/bri_timer_0/count_n2 , 
        \PLUSE_0/bri_coder_0/un2lto7_3_net_1 , 
        \PLUSE_0/bri_coder_0/un2lto7_1_net_1 , 
        \PLUSE_0/bri_coder_0/un2lto7_2_net_1 , 
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[1] , 
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[2] , 
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[0] , 
        \PLUSE_0/bri_coder_0/N_11 , \PLUSE_0/bri_coder_0/N_10 , 
        \PLUSE_0/bri_coder_0/N_9 , \PLUSE_0/bri_coder_0/N_6 , 
        \PLUSE_0/bri_coder_0/N_8 , \PLUSE_0/bri_coder_0/N_7 , 
        \PLUSE_0/bri_coder_0/N_5 , \PLUSE_0/bri_coder_0/N_2 , 
        \PLUSE_0/bri_coder_0/N_3 , \PLUSE_0/bri_coder_0/N_4 , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[3] , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[4] , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[5] , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[0] , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[1] , 
        \PLUSE_0/bri_coder_0/ACT_LT3_E[2] , 
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[2] , 
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[1] , 
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[0] , 
        \PLUSE_0/qq_state_1/stateover_0_sqmuxa_i_0 , 
        \PLUSE_0/qq_state_1/cs[3]_net_1 , 
        \PLUSE_0/qq_state_1/cs[4]_net_1 , 
        \PLUSE_0/qq_state_1/Q1Q8_Q2Q7_RNO_0_net_1 , 
        \PLUSE_0/qq_state_1/cs4 , \PLUSE_0/qq_state_1/cs_RNO_2[3] , 
        \PLUSE_0/qq_state_1/N_86 , \PLUSE_0/qq_state_1/N_87 , 
        \PLUSE_0/qq_state_1/cs_RNO_2[2] , \PLUSE_0/qq_state_1/N_89 , 
        \PLUSE_0/qq_state_1/N_88 , \PLUSE_0/qq_state_1/N_84 , 
        \PLUSE_0/qq_state_1/cs[1]_net_1 , 
        \PLUSE_0/qq_state_1/cs_RNO_2[1] , 
        \PLUSE_0/qq_state_1/cs_i[0]_net_1 , \PLUSE_0/qq_state_1/N_82 , 
        \PLUSE_0/qq_state_1/cs_RNO_3[4] , 
        \PLUSE_0/qq_state_1/stateover_RNO_1 , 
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 , 
        \PLUSE_0/qq_timer_0/count_n2 , \PLUSE_0/qq_timer_0/count_c1 , 
        \PLUSE_0/qq_timer_0/count_n3 , \PLUSE_0/qq_timer_0/count_c2 , 
        \PLUSE_0/qq_timer_0/count_n4 , \PLUSE_0/qq_timer_0/count_9_0 , 
        \PLUSE_0/qq_timer_0/count_n0 , \PLUSE_0/qq_timer_0/count_n1 , 
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 , 
        \PLUSE_0/qq_timer_1/count_n2 , \PLUSE_0/qq_timer_1/count_c1 , 
        \PLUSE_0/qq_timer_1/count_n3 , \PLUSE_0/qq_timer_1/count_c2 , 
        \PLUSE_0/qq_timer_1/count_n4 , \PLUSE_0/qq_timer_1/count_9_0 , 
        \PLUSE_0/qq_timer_1/count_n0 , \PLUSE_0/qq_timer_1/count_n1 , 
        \PLUSE_0/qq_coder_1/i_0_4[1] , \PLUSE_0/qq_coder_1/i_0_1[1] , 
        \PLUSE_0/qq_coder_1/i_0_2[1] , \PLUSE_0/qq_coder_1/i_0_0[1] , 
        \PLUSE_0/qq_coder_1/un1_count_1[0] , 
        \PLUSE_0/qq_coder_1/i_reg10_NE_3[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_2[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_3[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_NE_0[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_NE_2[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_0[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_2[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_0[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_1[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_2[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_0[0]_net_1 , 
        \PLUSE_0/qq_coder_1/i_reg10_NE[0]_net_1 , 
        \PLUSE_0/qq_coder_1/un1_qq_para2_i[0] , 
        \PLUSE_0/qq_coder_1/i_RNO_3[2] , 
        \PLUSE_0/qq_coder_1/i_RNO_7[1] , 
        \PLUSE_0/qq_coder_1/i_RNO_8[0] , 
        \PLUSE_0/qq_coder_1/i_RNO_3[3] , 
        \PLUSE_0/bri_state_0/csse_2_0_1 , \PLUSE_0/bri_state_0/N_144 , 
        \PLUSE_0/bri_state_0/csse_2_0_0 , 
        \PLUSE_0/bri_state_0/cs[3]_net_1 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_1_0 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_11 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_6 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_5 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_10 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_4 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_3 , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_7 , 
        \PLUSE_0/bri_state_0/cs[8]_net_1 , 
        \PLUSE_0/bri_state_0/cs[2]_net_1 , 
        \PLUSE_0/bri_state_0/cs_i_0[7] , 
        \PLUSE_0/bri_state_0/cs_i_0[13] , 
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_1 , 
        \PLUSE_0/bri_state_0/cs[4]_net_1 , 
        \PLUSE_0/bri_state_0/cs[5]_net_1 , 
        \PLUSE_0/bri_state_0/cs[9]_net_1 , 
        \PLUSE_0/bri_state_0/cs_i_0[12] , 
        \PLUSE_0/bri_state_0/cs_i_0[6] , \PLUSE_0/bri_state_0/N_181 , 
        \PLUSE_0/bri_state_0/csse_10_0_a4_0_0 , 
        \PLUSE_0/bri_state_0/cs[10]_net_1 , 
        \PLUSE_0/bri_state_0/N_142 , 
        \PLUSE_0/bri_state_0/csse_4_0_a4_0_0 , 
        \PLUSE_0/bri_state_0/cs[1]_net_1 , 
        \PLUSE_0/bri_state_0/csse_1_0_a4_0_0 , 
        \PLUSE_0/bri_state_0/cs[0]_net_1 , 
        \PLUSE_0/bri_state_0/cs_ns_e[3] , \PLUSE_0/bri_state_0/N_183 , 
        \PLUSE_0/bri_state_0/down30 , \PLUSE_0/bri_state_0/N_178 , 
        \PLUSE_0/bri_state_0/N_145 , \PLUSE_0/bri_state_0/N_180 , 
        \PLUSE_0/bri_state_0/csse_0_0_0_tz , 
        \PLUSE_0/bri_state_0/cs_ns_e[1] , 
        \PLUSE_0/bri_state_0/en_net_1 , 
        \PLUSE_0/bri_state_0/cs_ns_e[0] , \PLUSE_0/bri_state_0/N_179 , 
        \PLUSE_0/bri_state_0/cs[11]_net_1 , 
        \PLUSE_0/bri_state_0/cs_RNO[14]_net_1 , 
        \PLUSE_0/bri_state_0/cs[14]_net_1 , 
        \PLUSE_0/bri_state_0/cs_RNO[13]_net_1 , 
        \PLUSE_0/bri_state_0/cs_RNO_0[12] , 
        \PLUSE_0/bri_state_0/cs_ns_e[11] , 
        \PLUSE_0/bri_state_0/cs_RNO_0[10] , 
        \PLUSE_0/bri_state_0/cs_ns_e[9] , 
        \PLUSE_0/bri_state_0/cs_RNO_1[8] , 
        \PLUSE_0/bri_state_0/cs_RNO_0[7] , 
        \PLUSE_0/bri_state_0/cs_RNO_1[6] , 
        \PLUSE_0/bri_state_0/down32 , \PLUSE_0/bri_state_0/cs_ns_e[2] , 
        \PLUSE_0/bri_state_0/cs_RNO_4[4] , 
        \PLUSE_0/bri_state_0/cs_ns_e[5] , 
        \state_1ms_0/timecount_8_iv_2[6] , 
        \state_1ms_0/S_DUMPTIME[6]_net_1 , \state_1ms_0/CS[7]_net_1 , 
        \state_1ms_0/CUTTIME_i_m[6] , 
        \state_1ms_0/timecount_8_iv_1[6] , 
        \state_1ms_0/PLUSECYCLE[6]_net_1 , \state_1ms_0/CS[4]_net_1 , 
        \state_1ms_0/PLUSETIME_i_m[6] , 
        \state_1ms_0/timecount_8_iv_0[6] , 
        \state_1ms_0/M_DUMPTIME[6]_net_1 , \state_1ms_0/CS[6]_net_1 , 
        \state_1ms_0/CS_i[0]_net_1 , \state_1ms_0/timecount_8_iv_2[5] , 
        \state_1ms_0/S_DUMPTIME[5]_net_1 , 
        \state_1ms_0/CUTTIME_i_m[5] , 
        \state_1ms_0/timecount_8_iv_1[5] , 
        \state_1ms_0/PLUSECYCLE[5]_net_1 , 
        \state_1ms_0/PLUSETIME_i_m[5] , 
        \state_1ms_0/timecount_8_iv_0[5] , 
        \state_1ms_0/M_DUMPTIME[5]_net_1 , 
        \state_1ms_0/timecount_8_iv_2[1] , 
        \state_1ms_0/S_DUMPTIME[1]_net_1 , \state_1ms_0/CUTTIME_m[1] , 
        \state_1ms_0/timecount_8_iv_1[1] , 
        \state_1ms_0/PLUSECYCLE[1]_net_1 , 
        \state_1ms_0/PLUSETIME_m[1] , 
        \state_1ms_0/timecount_8_iv_0[1] , 
        \state_1ms_0/M_DUMPTIME[1]_net_1 , 
        \state_1ms_0/timecount_8_iv_2[3] , 
        \state_1ms_0/S_DUMPTIME[3]_net_1 , \state_1ms_0/CUTTIME_m[3] , 
        \state_1ms_0/timecount_8_iv_1[3] , 
        \state_1ms_0/PLUSECYCLE[3]_net_1 , 
        \state_1ms_0/PLUSETIME_m[3] , 
        \state_1ms_0/timecount_8_iv_0[3] , 
        \state_1ms_0/M_DUMPTIME[3]_net_1 , 
        \state_1ms_0/timecount_8_iv_2[2] , 
        \state_1ms_0/S_DUMPTIME[2]_net_1 , 
        \state_1ms_0/CUTTIME_i_m[2] , 
        \state_1ms_0/timecount_8_iv_1[2] , 
        \state_1ms_0/PLUSECYCLE[2]_net_1 , 
        \state_1ms_0/PLUSETIME_i_m[2] , 
        \state_1ms_0/timecount_8_iv_0[2] , 
        \state_1ms_0/M_DUMPTIME[2]_net_1 , 
        \state_1ms_0/timecount_8_0_iv_1[15] , 
        \state_1ms_0/S_DUMPTIME[15]_net_1 , 
        \state_1ms_0/PLUSETIME_m[15] , 
        \state_1ms_0/timecount_8_0_iv_0[15] , 
        \state_1ms_0/M_DUMPTIME[15]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[15] , 
        \state_1ms_0/timecount_8_0_iv_1[9] , 
        \state_1ms_0/S_DUMPTIME[9]_net_1 , 
        \state_1ms_0/PLUSETIME_m[9] , 
        \state_1ms_0/timecount_8_0_iv_0[9] , 
        \state_1ms_0/M_DUMPTIME[9]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[9] , 
        \state_1ms_0/timecount_8_0_iv_1[14] , 
        \state_1ms_0/S_DUMPTIME[14]_net_1 , 
        \state_1ms_0/PLUSETIME_m[14] , 
        \state_1ms_0/timecount_8_0_iv_0[14] , 
        \state_1ms_0/M_DUMPTIME[14]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[14] , 
        \state_1ms_0/timecount_8_0_iv_1[7] , 
        \state_1ms_0/S_DUMPTIME[7]_net_1 , 
        \state_1ms_0/PLUSETIME_m[7] , 
        \state_1ms_0/timecount_8_0_iv_0[7] , 
        \state_1ms_0/M_DUMPTIME[7]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[7] , 
        \state_1ms_0/timecount_8_0_iv_1[10] , 
        \state_1ms_0/S_DUMPTIME[10]_net_1 , 
        \state_1ms_0/PLUSETIME_m[10] , 
        \state_1ms_0/timecount_8_0_iv_0[10] , 
        \state_1ms_0/M_DUMPTIME[10]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[10] , 
        \state_1ms_0/timecount_8_0_iv_1[12] , 
        \state_1ms_0/S_DUMPTIME[12]_net_1 , 
        \state_1ms_0/PLUSETIME_m[12] , 
        \state_1ms_0/timecount_8_0_iv_0[12] , 
        \state_1ms_0/M_DUMPTIME[12]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[12] , 
        \state_1ms_0/timecount_8_0_iv_1[11] , 
        \state_1ms_0/S_DUMPTIME[11]_net_1 , 
        \state_1ms_0/PLUSETIME_m[11] , 
        \state_1ms_0/timecount_8_0_iv_0[11] , 
        \state_1ms_0/M_DUMPTIME[11]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[11] , 
        \state_1ms_0/timecount_8_0_iv_1[4] , 
        \state_1ms_0/S_DUMPTIME[4]_net_1 , 
        \state_1ms_0/PLUSETIME_m[4] , 
        \state_1ms_0/timecount_8_0_iv_0[4] , 
        \state_1ms_0/M_DUMPTIME[4]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[4] , 
        \state_1ms_0/timecount_8_0_iv_1[13] , 
        \state_1ms_0/S_DUMPTIME[13]_net_1 , 
        \state_1ms_0/PLUSETIME_m[13] , 
        \state_1ms_0/timecount_8_0_iv_0[13] , 
        \state_1ms_0/M_DUMPTIME[13]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[13] , 
        \state_1ms_0/timecount_8_0_iv_1[0] , 
        \state_1ms_0/S_DUMPTIME[0]_net_1 , 
        \state_1ms_0/PLUSETIME_m[0] , 
        \state_1ms_0/timecount_8_0_iv_0[0] , 
        \state_1ms_0/M_DUMPTIME[0]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[0] , 
        \state_1ms_0/timecount_8_0_iv_1[8] , 
        \state_1ms_0/S_DUMPTIME[8]_net_1 , 
        \state_1ms_0/PLUSETIME_m[8] , 
        \state_1ms_0/timecount_8_0_iv_0[8] , 
        \state_1ms_0/M_DUMPTIME[8]_net_1 , 
        \state_1ms_0/PLUSECYCLE_m[8] , \state_1ms_0/CS_srsts_i_0[9] , 
        \state_1ms_0/CS[8]_net_1 , \state_1ms_0/CS_srsts_i_0[8] , 
        \state_1ms_0/CS_srsts_i_0[1] , \state_1ms_0/CS_srsts_i_0[2] , 
        \state_1ms_0/CS[1]_net_1 , \state_1ms_0/CS_srsts_i_0[5] , 
        \state_1ms_0/CS_srsts_i_0[4] , \state_1ms_0/CS[3]_net_1 , 
        \state_1ms_0/CS_srsts_i_0[3] , \state_1ms_0/CS[2]_net_1 , 
        \state_1ms_0/CS_srsts_i_0[7] , \state_1ms_0/N_204s_i_i_0 , 
        \state_1ms_0/CS_srsts_i_0[6] , \state_1ms_0/CS[5]_net_1 , 
        \state_1ms_0/un1_CS_9_0_a4_0 , 
        \state_1ms_0/un1_PLUSECYCLE13_i_a2_0_net_1 , 
        \state_1ms_0/timecount_8[3] , \state_1ms_0/timecount_8_iv[2] , 
        \state_1ms_0/N_256 , \state_1ms_0/timecount_8[9] , 
        \state_1ms_0/CUTTIME_m[9] , \state_1ms_0/timecount_8[7] , 
        \state_1ms_0/CUTTIME_m[7] , \state_1ms_0/CS_RNO_1[8] , 
        \state_1ms_0/CS_RNO_3[1] , \state_1ms_0/CS_RNO_3[4] , 
        \state_1ms_0/CS_RNO_3[3] , \state_1ms_0/CS_RNO_3[2] , 
        \state_1ms_0/CS_RNO_3[5] , \state_1ms_0/CS_RNO_1[9] , 
        \state_1ms_0/CS[9]_net_1 , \state_1ms_0/CS_RNO_3[6] , 
        \state_1ms_0/CS_RNO_3[7] , \state_1ms_0/CS_i_RNO_1[0] , 
        \state_1ms_0/S_DUMPTIME_1_sqmuxa , \state_1ms_0/N_17 , 
        \state_1ms_0/PLUSETIME_1_sqmuxa , 
        \state_1ms_0/PLUSECYCLE_0_sqmuxa , 
        \state_1ms_0/M_DUMPTIME_1_sqmuxa , 
        \state_1ms_0/timecount_8[4] , \state_1ms_0/CUTTIME_m[4] , 
        \state_1ms_0/timecount_8[0] , \state_1ms_0/CUTTIME_m[0] , 
        \state_1ms_0/timecount_8[1] , \state_1ms_0/timecount_8_iv[5] , 
        \state_1ms_0/timecount_8_iv[6] , \state_1ms_0/timecount_8[10] , 
        \state_1ms_0/CUTTIME_m[10] , \state_1ms_0/timecount_8[14] , 
        \state_1ms_0/CUTTIME_m[14] , \state_1ms_0/timecount_8[8] , 
        \state_1ms_0/CUTTIME_m[8] , \state_1ms_0/timecount_8[11] , 
        \state_1ms_0/CUTTIME_m[11] , \state_1ms_0/timecount_8[12] , 
        \state_1ms_0/CUTTIME_m[12] , \state_1ms_0/timecount_8[13] , 
        \state_1ms_0/CUTTIME_m[13] , \state_1ms_0/timecount_8[15] , 
        \state_1ms_0/CUTTIME_m[15] , \state_1ms_0/N_154 , 
        \state_1ms_0/N_257 , \state_1ms_0/N_155 , \state_1ms_0/N_254 , 
        \state_1ms_0/N_156 , \state_1ms_0/bri_cycle_RNO_0_net_1 , 
        \state_1ms_0/pluse_start_RNO_2 , \state_1ms_0/reset_out_RNO_1 , 
        \state_1ms_0/timecount_RNO[1]_net_1 , \state_1ms_0/N_68 , 
        \state_1ms_0/timecount_RNO[4]_net_1 , \state_1ms_0/N_71 , 
        \state_1ms_0/timecount_RNO[5]_net_1 , \state_1ms_0/N_72 , 
        \state_1ms_0/timecount_RNO[6]_net_1 , \state_1ms_0/N_73 , 
        \state_1ms_0/timecount_RNO[8]_net_1 , \state_1ms_0/N_75 , 
        \state_1ms_0/timecount_RNO[10]_net_1 , \state_1ms_0/N_77 , 
        \state_1ms_0/timecount_RNO[11]_net_1 , \state_1ms_0/N_78 , 
        \state_1ms_0/timecount_RNO[12]_net_1 , \state_1ms_0/N_79 , 
        \state_1ms_0/timecount_RNO[13]_net_1 , \state_1ms_0/N_80 , 
        \state_1ms_0/timecount_RNO[14]_net_1 , \state_1ms_0/N_81 , 
        \state_1ms_0/timecount_RNO[15]_net_1 , \state_1ms_0/N_82 , 
        \state_1ms_0/timecount_RNO[0]_net_1 , \state_1ms_0/N_67 , 
        \state_1ms_0/N_16 , \state_1ms_0/PLUSECYCLE[8]_net_1 , 
        \state_1ms_0/PLUSETIME[8]_net_1 , 
        \state_1ms_0/CUTTIME[8]_net_1 , 
        \state_1ms_0/PLUSECYCLE[11]_net_1 , 
        \state_1ms_0/PLUSETIME[11]_net_1 , 
        \state_1ms_0/CUTTIME[11]_net_1 , 
        \state_1ms_0/PLUSECYCLE[12]_net_1 , 
        \state_1ms_0/PLUSETIME[12]_net_1 , 
        \state_1ms_0/CUTTIME[12]_net_1 , 
        \state_1ms_0/PLUSECYCLE[13]_net_1 , 
        \state_1ms_0/PLUSETIME[13]_net_1 , 
        \state_1ms_0/CUTTIME[13]_net_1 , 
        \state_1ms_0/PLUSECYCLE[15]_net_1 , 
        \state_1ms_0/PLUSETIME[15]_net_1 , 
        \state_1ms_0/CUTTIME[15]_net_1 , 
        \state_1ms_0/PLUSECYCLE[0]_net_1 , 
        \state_1ms_0/PLUSETIME[0]_net_1 , 
        \state_1ms_0/CUTTIME[0]_net_1 , 
        \state_1ms_0/PLUSETIME[1]_net_1 , 
        \state_1ms_0/CUTTIME[1]_net_1 , 
        \state_1ms_0/PLUSETIME[5]_net_1 , 
        \state_1ms_0/CUTTIME[5]_net_1 , 
        \state_1ms_0/PLUSETIME[6]_net_1 , 
        \state_1ms_0/CUTTIME[6]_net_1 , 
        \state_1ms_0/PLUSECYCLE[10]_net_1 , 
        \state_1ms_0/PLUSETIME[10]_net_1 , 
        \state_1ms_0/CUTTIME[10]_net_1 , 
        \state_1ms_0/PLUSECYCLE[14]_net_1 , 
        \state_1ms_0/PLUSETIME[14]_net_1 , 
        \state_1ms_0/CUTTIME[14]_net_1 , 
        \state_1ms_0/CUTTIME[4]_net_1 , 
        \state_1ms_0/PLUSETIME[4]_net_1 , 
        \state_1ms_0/PLUSECYCLE[4]_net_1 , \state_1ms_0/N_364 , 
        \state_1ms_0/N_380 , \state_1ms_0/N_255 , 
        \state_1ms_0/CUTTIME[9]_net_1 , 
        \state_1ms_0/PLUSETIME[9]_net_1 , 
        \state_1ms_0/PLUSECYCLE[9]_net_1 , 
        \state_1ms_0/CUTTIME[7]_net_1 , 
        \state_1ms_0/PLUSETIME[7]_net_1 , 
        \state_1ms_0/PLUSECYCLE[7]_net_1 , 
        \state_1ms_0/timecount_8[17] , \state_1ms_0/CUTTIME[17]_net_1 , 
        \state_1ms_0/timecount_8[19] , \state_1ms_0/CUTTIME[19]_net_1 , 
        \state_1ms_0/timecount_8[18] , \state_1ms_0/CUTTIME[18]_net_1 , 
        \state_1ms_0/timecount_8[16] , \state_1ms_0/CUTTIME[16]_net_1 , 
        \state_1ms_0/N_86 , \state_1ms_0/N_85 , \state_1ms_0/N_84 , 
        \state_1ms_0/N_83 , \state_1ms_0/N_76 , \state_1ms_0/N_74 , 
        \state_1ms_0/timecount_RNO[19]_net_1 , 
        \state_1ms_0/timecount_RNO[18]_net_1 , 
        \state_1ms_0/timecount_RNO[17]_net_1 , 
        \state_1ms_0/timecount_RNO[16]_net_1 , 
        \state_1ms_0/timecount_RNO[9]_net_1 , 
        \state_1ms_0/timecount_RNO[7]_net_1 , 
        \state_1ms_0/dump_start_RNO_2_net_1 , \state_1ms_0/N_87 , 
        \state_1ms_0/soft_dump_RNO_net_1 , \state_1ms_0/N_152 , 
        \state_1ms_0/rt_sw_RNO_3 , \state_1ms_0/N_153 , 
        \state_1ms_0/CUTTIME[3]_net_1 , 
        \state_1ms_0/PLUSETIME[3]_net_1 , 
        \state_1ms_0/CUTTIME[2]_net_1 , 
        \state_1ms_0/PLUSETIME[2]_net_1 , \state_1ms_0/N_70 , 
        \state_1ms_0/N_69 , \state_1ms_0/timecount_RNO[3]_net_1 , 
        \state_1ms_0/timecount_RNO[2]_net_1 , \sd_acq_top_0/i[9] , 
        \sd_acq_top_0/i[10] , \sd_acq_top_0/i_0[6] , 
        \sd_acq_top_0/i_0[7] , \sd_acq_top_0/i_0[8] , 
        \sd_acq_top_0/i_1[5] , \sd_acq_top_0/i_2[4] , 
        \sd_acq_top_0/i_5[2] , \sd_acq_top_0/i_5[3] , 
        \sd_acq_top_0/i_10[0] , \sd_acq_top_0/count[16] , 
        \sd_acq_top_0/count[17] , \sd_acq_top_0/count[18] , 
        \sd_acq_top_0/count[19] , \sd_acq_top_0/count[20] , 
        \sd_acq_top_0/count[21] , \sd_acq_top_0/count_0[12] , 
        \sd_acq_top_0/count_0[13] , \sd_acq_top_0/count_0[14] , 
        \sd_acq_top_0/count_0[15] , \sd_acq_top_0/count_1[8] , 
        \sd_acq_top_0/count_1[9] , \sd_acq_top_0/count_1[10] , 
        \sd_acq_top_0/count_1[11] , \sd_acq_top_0/count_10[0] , 
        \sd_acq_top_0/count_10[1] , \sd_acq_top_0/count_10[2] , 
        \sd_acq_top_0/count_10[3] , \sd_acq_top_0/count_10[4] , 
        \sd_acq_top_0/count_3[5] , \sd_acq_top_0/count_3[6] , 
        \sd_acq_top_0/count_3[7] , 
        \sd_acq_top_0/sd_sacq_state_0_stateover , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_21[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_18[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_17[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_19[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_8[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_7[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_16[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_4[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_3[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_14[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_2[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_1[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_11[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_10[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_6[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[10] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_2[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[18]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_14[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[16]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_19[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[20]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[21]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[8] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[6] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_3_i_a2_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_14[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_2[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_12[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_2[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_16[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_22[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_22[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[16]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_14[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[20]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_19[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[21]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_19[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_12[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_16[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_16[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_0_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[20]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_19[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[21]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_2[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_16[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_0_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_10[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_15[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[16]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_18[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[20]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_19[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[21]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_17[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_14[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_14[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_12[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_13[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_12[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_1[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_7[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_2[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_3[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_0[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_6[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_12[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_4[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_5[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_11[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_8[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_2[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_1[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_0[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_1_i_a2_0_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_i_a2_0_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa , 
        \sd_acq_top_0/sd_sacq_coder_0/N_23 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[7] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa , 
        \sd_acq_top_0/sd_sacq_coder_0/N_24 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_i[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[5] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[2] , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[3] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[16]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[17]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[17]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[17]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[19]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[19]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[19]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[18]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[18]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[4] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[3]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_366 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_382 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_394 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_404 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_410 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_426 , 
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_9[0] , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa , 
        \sd_acq_top_0/sd_sacq_coder_0/N_360 , 
        \sd_acq_top_0/sd_sacq_coder_0/N_344 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[18]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[19]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[17]_net_1 , 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[12] , 
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs4 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[9] , 
        \sd_acq_top_0/sd_sacq_state_0/en2_0_0_o3_0 , 
        \sd_acq_top_0/sd_sacq_state_0/N_233 , 
        \sd_acq_top_0/sd_sacq_state_0/N_232 , 
        \sd_acq_top_0/sd_sacq_state_0/N_201 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[4]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[11]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/ns_0_1_i_a2_0 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[14]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/N_245 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[2] , 
        \sd_acq_top_0/sd_sacq_state_0/N_214 , 
        \sd_acq_top_0/sd_sacq_state_0/N_215 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_5[4] , 
        \sd_acq_top_0/sd_sacq_state_0/en1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[5] , 
        \sd_acq_top_0/sd_sacq_state_0/N_216 , 
        \sd_acq_top_0/sd_sacq_state_0/N_217 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[6] , 
        \sd_acq_top_0/sd_sacq_state_0/N_218 , 
        \sd_acq_top_0/sd_sacq_state_0/N_219 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[8] , 
        \sd_acq_top_0/sd_sacq_state_0/N_221 , 
        \sd_acq_top_0/sd_sacq_state_0/N_222 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/N_207 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[9]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[11] , 
        \sd_acq_top_0/sd_sacq_state_0/cs[10]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/N_208 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[12]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[14] , 
        \sd_acq_top_0/sd_sacq_state_0/cs[13]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[3] , 
        \sd_acq_top_0/sd_sacq_state_0/N_237 , 
        \sd_acq_top_0/sd_sacq_state_0/N_236 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[1] , 
        \sd_acq_top_0/sd_sacq_state_0/cs_i[0]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[2]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[1]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[6]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[7] , 
        \sd_acq_top_0/sd_sacq_state_0/N_203 , 
        \sd_acq_top_0/sd_sacq_state_0/cs[7]_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[10] , 
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[13] , 
        \sd_acq_top_0/sd_sacq_state_0/en2_RNO_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/N_230 , 
        \sd_acq_top_0/sd_sacq_state_0/N_235 , 
        \sd_acq_top_0/sd_sacq_state_0/en2_net_1 , 
        \sd_acq_top_0/sd_sacq_state_0/stateover_RNO_2 , 
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO[15]_net_1 , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[21] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[21] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[20] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[20] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[19] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[19] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[18] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[18] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[17] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[17] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[16] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[16] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[15] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[15] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[14] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[14] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[13] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[13] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[12] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[12] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[11] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[11] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[10] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[10] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[9] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[9] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[8] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[8] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[7] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[7] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[6] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[6] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[5] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[5] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[4] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[4] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[3] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[3] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[2] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[2] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[1] , 
        \sd_acq_top_0/sd_sacq_timer_0/count1[1] , 
        \sd_acq_top_0/sd_sacq_timer_0/count_3[0] , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_16_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_5_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_8_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_8_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_7_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_17_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc1_25_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_16_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_27_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_19_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_9_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_5_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_12_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_13_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_10_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_15_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_11_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_14_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_14_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_20_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_24_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_20_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_31_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_21_net , 
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_33_net , 
        \syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en , 
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_i , 
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_net_1 , 
        \syn_md_module_1/syn_md_edge_detect_0/sig_r1_i_0 , 
        \syn_md_module_1/syn_md_combine_0/syn_md_temp_0_net_1 , 
        \syn_md_module_1/syn_md_0/count_n2_i_0 , 
        \syn_md_module_1/syn_md_0/count_n2_i_a2_0 , 
        \syn_md_module_1/syn_md_0/N_23_1 , 
        \syn_md_module_1/syn_md_0/count[0]_net_1 , 
        \syn_md_module_1/syn_md_0/count[1]_net_1 , 
        \syn_md_module_1/syn_md_0/count[2]_net_1 , 
        \syn_md_module_1/syn_md_0/N_14 , 
        \syn_md_module_1/syn_md_0/N_30 , 
        \syn_md_module_1/syn_md_0/N_31 , 
        \syn_md_module_1/syn_md_0/count_RNO_0[1]_net_1 , 
        \syn_md_module_1/syn_md_0/N_52 , 
        \syn_md_module_1/syn_md_0/N_18 , 
        \syn_md_module_1/syn_md_0/N_50 , 
        \syn_md_module_1/syn_md_0/count[3]_net_1 , 
        \syn_md_module_1/syn_md_0/N_28 , 
        \syn_md_module_1/syn_md_0/N_25 , 
        \syn_md_module_1/syn_md_0/N_22 , 
        \syn_md_module_1/syn_md_0/count_RNO_0[0]_net_1 , 
        \syn_md_module_1/syn_md_0/count_RNO[1]_net_1 , 
        \syn_md_module_1/syn_md_0/count_RNO[2]_net_1 , 
        \syn_md_module_1/syn_md_0/count_RNO[3]_net_1 , 
        \DUMP_OFF_1/i_4[0] , \DUMP_OFF_1/i_4[1] , 
        \DUMP_OFF_1/off_on_state_0_state_over , 
        \DUMP_OFF_1/count_4[0] , \DUMP_OFF_1/count_4[1] , 
        \DUMP_OFF_1/count_4[2] , \DUMP_OFF_1/count_4[3] , 
        \DUMP_OFF_1/count_4[4] , \DUMP_OFF_1/off_on_state_0/N_36_i , 
        \DUMP_OFF_1/off_on_state_0/N_42_i , 
        \DUMP_OFF_1/off_on_state_0/cs_nsss[1] , 
        \DUMP_OFF_1/off_on_state_0/N_10 , 
        \DUMP_OFF_1/off_on_state_0/cs[1]_net_1 , 
        \DUMP_OFF_1/off_on_state_0/N_9 , 
        \DUMP_OFF_1/off_on_state_0/N_12_mux , 
        \DUMP_OFF_1/off_on_coder_0/i_0_2[1] , 
        \DUMP_OFF_1/off_on_coder_0/i_0_1[1] , 
        \DUMP_OFF_1/off_on_coder_0/i_RNO_4[1] , 
        \DUMP_OFF_1/off_on_coder_0/i_RNO_4[0] , 
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 , 
        \DUMP_OFF_1/off_on_timer_0/count_n2 , 
        \DUMP_OFF_1/off_on_timer_0/count_c1 , 
        \DUMP_OFF_1/off_on_timer_0/count_n3 , 
        \DUMP_OFF_1/off_on_timer_0/count_c2 , 
        \DUMP_OFF_1/off_on_timer_0/count_n4 , 
        \DUMP_OFF_1/off_on_timer_0/count_9_0 , 
        \DUMP_OFF_1/off_on_timer_0/count_n0 , 
        \DUMP_OFF_1/off_on_timer_0/count_n1 , 
        \scalestate_0/CS_0[11]_net_1 , 
        \scalestate_0/CS_RNIRUEO[10]_net_1 , 
        \scalestate_0/un1_CS6_33_2 , \scalestate_0/N_1310 , 
        \scalestate_0/un1_CS6_33_1 , \scalestate_0/un1_CS6_33_0 , 
        \scalestate_0/N_258_0 , \scalestate_0/timecount_12_sqmuxa_0 , 
        \scalestate_0/N_1209_0 , \scalestate_0/N_1194 , 
        \scalestate_0/N_1265 , 
        \scalestate_0/un1_timecount_2_sqmuxa_7_reto , 
        \scalestate_0/un1_timecount_2_sqmuxa_7 , 
        \scalestate_0/un1_CS6_33 , 
        \scalestate_0/timecount_m3_e_2_reto , 
        \scalestate_0/timecount_m3_e_2 , 
        \scalestate_0/timecount_m3_e_1_reto , 
        \scalestate_0/timecount_m3_e_1 , 
        \scalestate_0/timecount_11_sqmuxa_m_reto , 
        \scalestate_0/timecount_20_iv_6_reto[8] , 
        \scalestate_0/timecount_20_iv_6[8] , 
        \scalestate_0/timecount_20_iv_2_reto[8] , 
        \scalestate_0/timecount_20_iv_2[8] , 
        \scalestate_0/timecount_20_iv_3_reto[8] , 
        \scalestate_0/timecount_20_iv_3[8] , 
        \scalestate_0/timecount_20_iv_9_reto[8] , 
        \scalestate_0/timecount_20_iv_6_reto[10] , 
        \scalestate_0/timecount_20_iv_6[10] , 
        \scalestate_0/timecount_20_iv_2_reto[10] , 
        \scalestate_0/timecount_20_iv_2[10] , 
        \scalestate_0/timecount_20_iv_3_reto[10] , 
        \scalestate_0/timecount_20_iv_3[10] , 
        \scalestate_0/timecount_20_iv_9_reto[10] , 
        \scalestate_0/timecount_20_iv_6_reto[11] , 
        \scalestate_0/timecount_20_iv_6[11] , 
        \scalestate_0/timecount_20_iv_2_reto[11] , 
        \scalestate_0/timecount_20_iv_2[11] , 
        \scalestate_0/timecount_20_iv_3_reto[11] , 
        \scalestate_0/timecount_20_iv_3[11] , 
        \scalestate_0/timecount_20_iv_9_reto[11] , 
        \scalestate_0/timecount_20_iv_6_reto[4] , 
        \scalestate_0/timecount_20_iv_6[4] , 
        \scalestate_0/timecount_20_iv_2_reto[4] , 
        \scalestate_0/timecount_20_iv_2[4] , 
        \scalestate_0/timecount_20_iv_3_reto[4] , 
        \scalestate_0/timecount_20_iv_3[4] , 
        \scalestate_0/timecount_20_iv_9_reto[4] , 
        \scalestate_0/un1_timecount_2_sqmuxa_9_reto , 
        \scalestate_0/un1_timecount_2_sqmuxa_9 , 
        \scalestate_0/timecount_m1_e_2_2_reto , 
        \scalestate_0/timecount_m1_e_2_2 , 
        \scalestate_0/timecount_cnst_m_reto[1] , 
        \scalestate_0/timecount_20_iv_8_reto[6] , 
        \scalestate_0/timecount_20_iv_8[6] , 
        \scalestate_0/timecount_20_iv_9_reto[6] , 
        \scalestate_0/timecount_20_iv_9[6] , 
        \scalestate_0/timecount_20_iv_10_reto[6] , 
        \scalestate_0/timecount_20_iv_8_reto[5] , 
        \scalestate_0/timecount_20_iv_8[5]_net_1 , 
        \scalestate_0/timecount_20_iv_9_reto[5] , 
        \scalestate_0/timecount_20_iv_9[5] , 
        \scalestate_0/timecount_20_iv_8_reto[7] , 
        \scalestate_0/timecount_20_iv_8[7] , 
        \scalestate_0/timecount_20_iv_6_reto[7] , 
        \scalestate_0/timecount_20_iv_6[7] , 
        \scalestate_0/timecount_20_iv_7_reto[7] , 
        \scalestate_0/timecount_20_iv_7[7] , 
        \scalestate_0/timecount_20_iv_10_reto[7] , 
        \scalestate_0/timecount_20_iv_8_reto[15] , 
        \scalestate_0/timecount_20_iv_8[15] , 
        \scalestate_0/timecount_20_iv_6_reto[15] , 
        \scalestate_0/timecount_20_iv_6[15] , 
        \scalestate_0/timecount_20_iv_7_reto[15] , 
        \scalestate_0/timecount_20_iv_7[15] , 
        \scalestate_0/timecount_20_iv_8_reto[14] , 
        \scalestate_0/timecount_20_iv_8[14] , 
        \scalestate_0/timecount_20_iv_6_reto[14] , 
        \scalestate_0/timecount_20_iv_6[14] , 
        \scalestate_0/timecount_20_iv_7_reto[14] , 
        \scalestate_0/timecount_20_iv_7[14] , 
        \scalestate_0/timecount_20_iv_8_reto[13] , 
        \scalestate_0/timecount_20_iv_8[13] , 
        \scalestate_0/timecount_20_iv_6_reto[13] , 
        \scalestate_0/timecount_20_iv_6[13] , 
        \scalestate_0/timecount_20_iv_7_reto[13] , 
        \scalestate_0/timecount_20_iv_7[13] , 
        \scalestate_0/timecount_20_iv_8_reto[12] , 
        \scalestate_0/timecount_20_iv_8[12] , 
        \scalestate_0/timecount_20_iv_6_reto[12] , 
        \scalestate_0/timecount_20_iv_6[12] , 
        \scalestate_0/timecount_20_iv_7_reto[12] , 
        \scalestate_0/timecount_20_iv_7[12] , 
        \scalestate_0/timecount_20_iv_8_reto[0] , 
        \scalestate_0/timecount_20_iv_8[0] , 
        \scalestate_0/timecount_20_iv_6_reto[0] , 
        \scalestate_0/timecount_20_iv_6[0] , 
        \scalestate_0/timecount_20_iv_7_reto[0] , 
        \scalestate_0/timecount_20_iv_7[0] , 
        \scalestate_0/timecount_20_0_iv_4_reto[19] , 
        \scalestate_0/timecount_20_0_iv_4[19] , 
        \scalestate_0/OPENTIME_TEL_m_reto[19] , 
        \scalestate_0/OPENTIME_TEL_m[19] , 
        \scalestate_0/timecount_20_0_iv_0_reto[19] , 
        \scalestate_0/timecount_20_0_iv_0[19] , 
        \scalestate_0/timecount_20_0_iv_4_reto[18] , 
        \scalestate_0/timecount_20_0_iv_4[18] , 
        \scalestate_0/OPENTIME_TEL_m_reto[18] , 
        \scalestate_0/OPENTIME_TEL_m[18] , 
        \scalestate_0/timecount_20_0_iv_0_reto[18] , 
        \scalestate_0/timecount_20_0_iv_0[18] , 
        \scalestate_0/timecount_20_0_iv_4_reto[17] , 
        \scalestate_0/timecount_20_0_iv_4[17] , 
        \scalestate_0/OPENTIME_TEL_m_reto[17] , 
        \scalestate_0/OPENTIME_TEL_m[17] , 
        \scalestate_0/timecount_20_0_iv_0_reto[17] , 
        \scalestate_0/timecount_20_0_iv_0[17] , 
        \scalestate_0/timecount_20_0_iv_4_reto[16] , 
        \scalestate_0/timecount_20_0_iv_4[16] , 
        \scalestate_0/OPENTIME_TEL_m_reto[16] , 
        \scalestate_0/OPENTIME_TEL_m[16] , 
        \scalestate_0/timecount_20_0_iv_0_reto[16] , 
        \scalestate_0/timecount_20_0_iv_0[16] , 
        \scalestate_0/un1_timecount_2_sqmuxa_1_reto , 
        \scalestate_0/un1_timecount_2_sqmuxa_1 , 
        \scalestate_0/un1_timecount_2_sqmuxa_reto , 
        \scalestate_0/timecount_20_iv_8_reto[2] , 
        \scalestate_0/timecount_20_iv_8[2] , 
        \scalestate_0/timecount_20_iv_6_reto[2] , 
        \scalestate_0/timecount_20_iv_6[2] , 
        \scalestate_0/timecount_20_iv_7_reto[2] , 
        \scalestate_0/timecount_20_iv_7[2] , 
        \scalestate_0/timecount_20_iv_10_reto[2] , 
        \scalestate_0/timecount_20_iv_8_reto[3] , 
        \scalestate_0/timecount_20_iv_8[3] , 
        \scalestate_0/timecount_20_iv_6_reto[3] , 
        \scalestate_0/timecount_20_iv_6[3] , 
        \scalestate_0/timecount_20_iv_7_reto[3] , 
        \scalestate_0/timecount_20_iv_7[3] , 
        \scalestate_0/timecount_20_iv_10_reto[3] , 
        \scalestate_0/timecount_20_iv_8_reto[9] , 
        \scalestate_0/timecount_20_iv_8[9] , 
        \scalestate_0/timecount_20_iv_6_reto[9] , 
        \scalestate_0/timecount_20_iv_6[9] , 
        \scalestate_0/timecount_20_iv_7_reto[9] , 
        \scalestate_0/timecount_20_iv_7[9] , 
        \scalestate_0/timecount_20_iv_10_reto[9] , 
        \scalestate_0/timecount_20_iv_8_reto[4] , 
        \scalestate_0/timecount_20_iv_8[4]_net_1 , 
        \scalestate_0/timecount_20_iv_8_reto[1] , 
        \scalestate_0/timecount_20_iv_8[1] , 
        \scalestate_0/timecount_20_iv_9_reto[1] , 
        \scalestate_0/timecount_20_iv_9[1] , 
        \scalestate_0/timecount_20_iv_8_reto[11] , 
        \scalestate_0/timecount_20_iv_8[11]_net_1 , 
        \scalestate_0/timecount_20_iv_8_reto[10] , 
        \scalestate_0/timecount_20_iv_8[10] , 
        \scalestate_0/timecount_20_iv_8_reto[8] , 
        \scalestate_0/timecount_20_iv_8[8] , 
        \scalestate_0/timecount_cnst_reto[5] , 
        \scalestate_0/timecount_cnst[5] , 
        \scalestate_0/timecount_cnst_m_reto[5] , 
        \scalestate_0/timecount_cnst_m_0_reto[6] , 
        \scalestate_0/timecount_cnst_m_0[6] , 
        \scalestate_0/timecount_cnst_m_reto[6] , 
        \scalestate_0/timecount_cnst_m_0_reto[9] , 
        \scalestate_0/timecount_cnst_m_0[9] , 
        \scalestate_0/timecount_cnst_m_0_reto[7] , 
        \scalestate_0/timecount_cnst_m_0[7] , 
        \scalestate_0/timecount_cnst_m_0_reto[3] , 
        \scalestate_0/timecount_cnst_m_0[3] , 
        \scalestate_0/timecount_cnst_m_0_reto[2] , 
        \scalestate_0/timecount_cnst_m_0[2] , 
        \scalestate_0/timecount_20_iv_0[5] , 
        \scalestate_0/OPENTIME_TEL_m[5] , 
        \scalestate_0/timecount_20_iv_4[5]_net_1 , 
        \scalestate_0/CUTTIMEI90_m[5] , 
        \scalestate_0/timecount_20_iv_4[11]_net_1 , 
        \scalestate_0/timecount_20_iv_0[11] , 
        \scalestate_0/OPENTIME_TEL_m[11] , 
        \scalestate_0/CUTTIMEI90_m[11] , 
        \scalestate_0/timecount_20_iv_5[4]_net_1 , 
        \scalestate_0/timecount_20_iv_4[4]_net_1 , 
        \scalestate_0/timecount_20_iv_0[4] , 
        \scalestate_0/CUTTIME90_m[4] , 
        \scalestate_0/timecount_20_iv_3[6] , 
        \scalestate_0/timecount_20_iv_2[6] , 
        \scalestate_0/timecount_20_iv_6[6] , 
        \scalestate_0/timecount_20_iv_0[6] , 
        \scalestate_0/OPENTIME_TEL_m[6] , 
        \scalestate_0/timecount_20_iv_4[6] , \scalestate_0/N_1089 , 
        \scalestate_0/S_DUMPTIME[6]_net_1 , 
        \scalestate_0/timecount_20_iv_1[6] , 
        \scalestate_0/CUTTIMEI90[6]_net_1 , \scalestate_0/N_252 , 
        \scalestate_0/CUTTIME90_m[6] , 
        \scalestate_0/CUTTIME180_TEL[6]_net_1 , \scalestate_0/N_261 , 
        \scalestate_0/CUTTIME180_Tini_m[6] , 
        \scalestate_0/OPENTIME[6]_net_1 , \scalestate_0/N_259 , 
        \scalestate_0/CUTTIME180_m[6] , \scalestate_0/N_1093 , 
        \scalestate_0/DUMPTIME[6]_net_1 , 
        \scalestate_0/PLUSETIME90_m[6] , \scalestate_0/N_1065 , 
        \scalestate_0/ACQTIME[6]_net_1 , 
        \scalestate_0/PLUSETIME180_m[6] , 
        \scalestate_0/timecount_20_iv_0[2] , 
        \scalestate_0/OPENTIME_TEL_m[2] , 
        \scalestate_0/timecount_20_iv_4[2] , 
        \scalestate_0/CUTTIME180_TEL_m[2] , 
        \scalestate_0/CUTTIME180_Tini_m[2] , 
        \scalestate_0/timecount_20_iv_2[2] , 
        \scalestate_0/S_DUMPTIME[2]_net_1 , 
        \scalestate_0/timecount_20_iv_1[2] , \scalestate_0/N_1069 , 
        \scalestate_0/CUTTIME90[2]_net_1 , 
        \scalestate_0/CUTTIMEI90_m[2] , 
        \scalestate_0/CUTTIME180[2]_net_1 , \scalestate_0/N_263 , 
        \scalestate_0/OPENTIME_m[2] , \scalestate_0/DUMPTIME[2]_net_1 , 
        \scalestate_0/PLUSETIME90_m[2] , 
        \scalestate_0/ACQTIME[2]_net_1 , 
        \scalestate_0/PLUSETIME180_m[2] , 
        \scalestate_0/timecount_20_iv_0[7] , 
        \scalestate_0/OPENTIME_TEL_m[7] , 
        \scalestate_0/timecount_20_iv_4[7] , 
        \scalestate_0/CUTTIME180_TEL_m[7] , 
        \scalestate_0/CUTTIME180_Tini_m[7] , 
        \scalestate_0/timecount_20_iv_2[7] , 
        \scalestate_0/S_DUMPTIME[7]_net_1 , 
        \scalestate_0/timecount_20_iv_1[7] , 
        \scalestate_0/CUTTIMEI90[7]_net_1 , 
        \scalestate_0/CUTTIME90_m[7] , 
        \scalestate_0/CUTTIME180[7]_net_1 , 
        \scalestate_0/OPENTIME_m[7] , \scalestate_0/DUMPTIME[7]_net_1 , 
        \scalestate_0/PLUSETIME90_m[7] , 
        \scalestate_0/ACQTIME[7]_net_1 , 
        \scalestate_0/PLUSETIME180_m[7] , 
        \scalestate_0/timecount_20_iv_0[3] , 
        \scalestate_0/OPENTIME_TEL_m[3] , 
        \scalestate_0/timecount_20_iv_4[3] , 
        \scalestate_0/CUTTIME180_TEL_m[3] , 
        \scalestate_0/CUTTIME180_Tini_m[3] , 
        \scalestate_0/timecount_20_iv_2[3] , 
        \scalestate_0/S_DUMPTIME[3]_net_1 , 
        \scalestate_0/timecount_20_iv_1[3] , 
        \scalestate_0/CUTTIME90[3]_net_1 , 
        \scalestate_0/CUTTIMEI90_m[3] , 
        \scalestate_0/CUTTIME180[3]_net_1 , 
        \scalestate_0/OPENTIME_m[3] , \scalestate_0/DUMPTIME[3]_net_1 , 
        \scalestate_0/PLUSETIME90_m[3] , 
        \scalestate_0/ACQTIME[3]_net_1 , 
        \scalestate_0/PLUSETIME180_m[3] , 
        \scalestate_0/CUTTIMEI90_m[9] , \scalestate_0/CUTTIME90_m[9] , 
        \scalestate_0/timecount_20_iv_5[9] , 
        \scalestate_0/CUTTIME180_TEL_m[9] , 
        \scalestate_0/CUTTIME180_Tini_m[9] , 
        \scalestate_0/timecount_20_iv_2[9] , 
        \scalestate_0/S_DUMPTIME[9]_net_1 , 
        \scalestate_0/timecount_20_iv_1[9] , 
        \scalestate_0/PLUSETIME180_m[9] , \scalestate_0/ACQTIME_m[9] , 
        \scalestate_0/OPENTIME_TEL_m[9] , 
        \scalestate_0/CUTTIME180[9]_net_1 , 
        \scalestate_0/OPENTIME_m[9] , \scalestate_0/DUMPTIME[9]_net_1 , 
        \scalestate_0/PLUSETIME90_m[9] , 
        \scalestate_0/timecount_20_iv_3[5] , 
        \scalestate_0/timecount_20_iv_2[5] , 
        \scalestate_0/timecount_20_iv_6[5] , 
        \scalestate_0/S_DUMPTIME[5]_net_1 , 
        \scalestate_0/timecount_20_iv_1[5] , 
        \scalestate_0/CUTTIME180_TEL[5]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[5] , 
        \scalestate_0/CUTTIME180[5]_net_1 , 
        \scalestate_0/OPENTIME_m[5] , \scalestate_0/DUMPTIME[5]_net_1 , 
        \scalestate_0/PLUSETIME90_m[5] , 
        \scalestate_0/ACQTIME[5]_net_1 , 
        \scalestate_0/PLUSETIME180_m[5] , \scalestate_0/N_1267 , 
        \scalestate_0/N_1197 , \scalestate_0/N_1206 , 
        \scalestate_0/un1_CS_20 , \scalestate_0/CS[16]_net_1 , 
        \scalestate_0/N_1153_1 , \scalestate_0/N_508_i_0_0 , 
        \scalestate_0/PLUSETIME90_m[11] , 
        \scalestate_0/DUMPTIME_m[11] , \scalestate_0/S_DUMPTIME_m[11] , 
        \scalestate_0/CUTTIME180_TEL[11]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[11] , 
        \scalestate_0/OPENTIME[11]_net_1 , 
        \scalestate_0/CUTTIME180_m[11] , 
        \scalestate_0/ACQTIME[11]_net_1 , 
        \scalestate_0/PLUSETIME180_m[11] , 
        \scalestate_0/timecount_20_iv_0[8] , 
        \scalestate_0/OPENTIME_TEL_m[8] , 
        \scalestate_0/timecount_20_iv_4[8] , 
        \scalestate_0/PLUSETIME90_m[8] , \scalestate_0/DUMPTIME_m[8] , 
        \scalestate_0/S_DUMPTIME_m[8] , 
        \scalestate_0/CUTTIMEI90[8]_net_1 , 
        \scalestate_0/CUTTIME90_m[8] , 
        \scalestate_0/CUTTIME180_TEL[8]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[8] , 
        \scalestate_0/CUTTIME180[8]_net_1 , 
        \scalestate_0/OPENTIME_m[8] , \scalestate_0/ACQTIME[8]_net_1 , 
        \scalestate_0/PLUSETIME180_m[8] , 
        \scalestate_0/timecount_20_iv_0[10] , 
        \scalestate_0/OPENTIME_TEL_m[10] , 
        \scalestate_0/timecount_20_iv_4[10] , 
        \scalestate_0/PLUSETIME90_m[10] , 
        \scalestate_0/DUMPTIME_m[10] , \scalestate_0/S_DUMPTIME_m[10] , 
        \scalestate_0/CUTTIMEI90[10]_net_1 , 
        \scalestate_0/CUTTIME90_m[10] , 
        \scalestate_0/CUTTIME180_TEL[10]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[10] , 
        \scalestate_0/OPENTIME[10]_net_1 , 
        \scalestate_0/CUTTIME180_m[10] , 
        \scalestate_0/ACQTIME[10]_net_1 , 
        \scalestate_0/PLUSETIME180_m[10] , 
        \scalestate_0/PLUSETIME90_m[4] , \scalestate_0/DUMPTIME_m[4] , 
        \scalestate_0/S_DUMPTIME_m[4] , 
        \scalestate_0/CUTTIME180_TEL[4]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[4] , 
        \scalestate_0/CUTTIME180[4]_net_1 , 
        \scalestate_0/OPENTIME_m[4] , \scalestate_0/ACQTIME[4]_net_1 , 
        \scalestate_0/PLUSETIME180_m[4] , 
        \scalestate_0/S_DUMPTIME_m[1] , 
        \scalestate_0/timecount_20_iv_1[1] , 
        \scalestate_0/timecount_20_iv_7[1] , 
        \scalestate_0/timecount_20_iv_0[1] , 
        \scalestate_0/OPENTIME_TEL_m[1] , 
        \scalestate_0/timecount_20_iv_4[1] , 
        \scalestate_0/OPENTIME_m[1] , \scalestate_0/CUTTIME180_m[1] , 
        \scalestate_0/timecount_20_iv_3[1] , 
        \scalestate_0/CUTTIMEI90[1]_net_1 , 
        \scalestate_0/CUTTIME90_m[1] , 
        \scalestate_0/CUTTIME180_TEL[1]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[1] , 
        \scalestate_0/DUMPTIME[1]_net_1 , 
        \scalestate_0/PLUSETIME90_m[1] , 
        \scalestate_0/ACQTIME[1]_net_1 , 
        \scalestate_0/PLUSETIME180_m[1] , 
        \scalestate_0/un1_timecount_2_sqmuxa_4 , 
        \scalestate_0/un1_timecount_2_sqmuxa_6_0 , 
        \scalestate_0/un1_timecount_2_sqmuxa_6_1 , 
        \scalestate_0/timecount_11_sqmuxa , 
        \scalestate_0/un1_CS6_26_0 , \scalestate_0/N_1209 , 
        \scalestate_0/fst_lst_pulse_net_1 , \scalestate_0/N_1196 , 
        \scalestate_0/timecount_m1_e_2_0 , 
        \scalestate_0/timecount_cnst[1] , 
        \scalestate_0/timecount_20_iv_0[12] , 
        \scalestate_0/OPENTIME_TEL_m[12] , 
        \scalestate_0/timecount_20_iv_4[12] , 
        \scalestate_0/CUTTIME180_m[12] , \scalestate_0/OPENTIME_m[12] , 
        \scalestate_0/timecount_20_iv_3[12] , 
        \scalestate_0/ACQTIME_m[12] , \scalestate_0/PLUSETIME90_m[12] , 
        \scalestate_0/S_DUMPTIME_m[12] , 
        \scalestate_0/CUTTIMEI90[12]_net_1 , 
        \scalestate_0/CUTTIME90_m[12] , 
        \scalestate_0/CUTTIME180_TEL[12]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[12] , 
        \scalestate_0/DUMPTIME[12]_net_1 , 
        \scalestate_0/PLUSETIME180_m[12] , 
        \scalestate_0/timecount_20_iv_0[13] , 
        \scalestate_0/OPENTIME_TEL_m[13] , 
        \scalestate_0/timecount_20_iv_4[13] , 
        \scalestate_0/CUTTIME180_m[13] , \scalestate_0/OPENTIME_m[13] , 
        \scalestate_0/timecount_20_iv_3[13] , 
        \scalestate_0/ACQTIME_m[13] , \scalestate_0/PLUSETIME90_m[13] , 
        \scalestate_0/S_DUMPTIME_m[13] , 
        \scalestate_0/CUTTIMEI90[13]_net_1 , 
        \scalestate_0/CUTTIME90_m[13] , 
        \scalestate_0/CUTTIME180_TEL[13]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[13] , 
        \scalestate_0/DUMPTIME[13]_net_1 , 
        \scalestate_0/PLUSETIME180_m[13] , 
        \scalestate_0/timecount_20_iv_0[0] , 
        \scalestate_0/OPENTIME_TEL_m[0] , 
        \scalestate_0/timecount_20_iv_4[0] , 
        \scalestate_0/CUTTIME180_m[0] , \scalestate_0/OPENTIME_m[0] , 
        \scalestate_0/timecount_20_iv_3[0] , 
        \scalestate_0/ACQTIME_m[0] , \scalestate_0/PLUSETIME90_m[0] , 
        \scalestate_0/S_DUMPTIME_m[0] , 
        \scalestate_0/CUTTIMEI90[0]_net_1 , 
        \scalestate_0/CUTTIME90_m[0] , 
        \scalestate_0/CUTTIME180_TEL[0]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[0] , 
        \scalestate_0/DUMPTIME[0]_net_1 , 
        \scalestate_0/PLUSETIME180_m[0] , 
        \scalestate_0/timecount_20_iv_0[14] , 
        \scalestate_0/OPENTIME_TEL_m[14] , 
        \scalestate_0/timecount_20_iv_4[14] , 
        \scalestate_0/CUTTIME180_m[14] , \scalestate_0/OPENTIME_m[14] , 
        \scalestate_0/timecount_20_iv_3[14] , 
        \scalestate_0/ACQTIME_m[14] , \scalestate_0/PLUSETIME90_m[14] , 
        \scalestate_0/S_DUMPTIME_m[14] , 
        \scalestate_0/CUTTIMEI90[14]_net_1 , 
        \scalestate_0/CUTTIME90_m[14] , 
        \scalestate_0/CUTTIME180_TEL[14]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[14] , 
        \scalestate_0/DUMPTIME[14]_net_1 , 
        \scalestate_0/PLUSETIME180_m[14] , 
        \scalestate_0/timecount_20_iv_0[15] , 
        \scalestate_0/OPENTIME_TEL_m[15] , 
        \scalestate_0/timecount_20_iv_4[15] , 
        \scalestate_0/CUTTIME180_m[15] , \scalestate_0/OPENTIME_m[15] , 
        \scalestate_0/timecount_20_iv_3[15] , 
        \scalestate_0/S_DUMPTIME[15]_net_1 , 
        \scalestate_0/timecount_20_iv_1[15] , 
        \scalestate_0/CUTTIMEI90[15]_net_1 , 
        \scalestate_0/CUTTIME90_m[15] , 
        \scalestate_0/CUTTIME180_TEL[15]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[15] , 
        \scalestate_0/ACQTIME[15]_net_1 , 
        \scalestate_0/PLUSETIME90_m[15] , 
        \scalestate_0/DUMPTIME[15]_net_1 , 
        \scalestate_0/PLUSETIME180_m[15] , 
        \scalestate_0/CUTTIME180_TEL_m[17] , 
        \scalestate_0/CUTTIME180_Tini_m[17] , 
        \scalestate_0/timecount_20_0_iv_2[17] , 
        \scalestate_0/CUTTIMEI90[17]_net_1 , 
        \scalestate_0/CUTTIME90_m[17] , 
        \scalestate_0/OPENTIME[17]_net_1 , 
        \scalestate_0/CUTTIME180_m[17] , 
        \scalestate_0/CUTTIME180_TEL_m[16] , 
        \scalestate_0/CUTTIME180_Tini_m[16] , 
        \scalestate_0/timecount_20_0_iv_2[16] , 
        \scalestate_0/CUTTIMEI90[16]_net_1 , 
        \scalestate_0/CUTTIME90_m[16] , 
        \scalestate_0/OPENTIME[16]_net_1 , 
        \scalestate_0/CUTTIME180_m[16] , 
        \scalestate_0/CUTTIME180_TEL_m[18] , 
        \scalestate_0/CUTTIME180_Tini_m[18] , 
        \scalestate_0/timecount_20_0_iv_2[18] , 
        \scalestate_0/CUTTIMEI90[18]_net_1 , 
        \scalestate_0/CUTTIME90_m[18] , 
        \scalestate_0/OPENTIME[18]_net_1 , 
        \scalestate_0/CUTTIME180_m[18] , 
        \scalestate_0/CUTTIME180_TEL_m[19] , 
        \scalestate_0/CUTTIME180_Tini_m[19] , 
        \scalestate_0/timecount_20_0_iv_2[19] , 
        \scalestate_0/CUTTIMEI90[19]_net_1 , 
        \scalestate_0/CUTTIME90_m[19] , 
        \scalestate_0/OPENTIME[19]_net_1 , 
        \scalestate_0/CUTTIME180_m[19] , 
        \scalestate_0/timecount_20_0_iv_1[21] , 
        \scalestate_0/CUTTIMEI90[21]_net_1 , 
        \scalestate_0/CUTTIME90_m[21] , 
        \scalestate_0/timecount_20_0_iv_0[21] , 
        \scalestate_0/CUTTIME180_TEL[21]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[21] , 
        \scalestate_0/timecount_20_0_iv_1[20] , 
        \scalestate_0/CUTTIMEI90[20]_net_1 , 
        \scalestate_0/CUTTIME90_m[20] , 
        \scalestate_0/timecount_20_0_iv_0[20] , 
        \scalestate_0/CUTTIME180_TEL[20]_net_1 , 
        \scalestate_0/CUTTIME180_Tini_m[20] , 
        \scalestate_0/un1_timecount_2_sqmuxa_7_0 , 
        \scalestate_0/necount_LE_M_RNIBQQD_net_1 , 
        \scalestate_0/CS[19]_net_1 , \scalestate_0/CS[14]_net_1 , 
        \scalestate_0/CS[20]_net_1 , 
        \scalestate_0/timecount_8_sqmuxa_i_0 , 
        \scalestate_0/CS[5]_net_1 , \scalestate_0/CS[13]_net_1 , 
        \scalestate_0/CS[12]_net_1 , \scalestate_0/necount_LE_M_net_1 , 
        \scalestate_0/timecount_17_sqmuxa_1 , 
        \scalestate_0/CS[15]_net_1 , \scalestate_0/M_pulse_net_1 , 
        \scalestate_0/timecount_13_sqmuxa_0 , 
        \scalestate_0/CS_srsts_i_0[8] , \scalestate_0/CS[8]_net_1 , 
        \scalestate_0/N_1263 , \scalestate_0/N_1210 , 
        \scalestate_0/un1_CS6_25_i_a3_0 , \scalestate_0/N_1266 , 
        \scalestate_0/N_1251_1 , \scalestate_0/CS_srsts_i_0[2] , 
        \scalestate_0/CS[2]_net_1 , \scalestate_0/N_1201 , 
        \scalestate_0/fst_lst_pulse8_NE_8 , 
        \scalestate_0/fst_lst_pulse8_NE_2 , 
        \scalestate_0/fst_lst_pulse8_NE_1 , 
        \scalestate_0/fst_lst_pulse8_NE_5 , 
        \scalestate_0/fst_lst_pulse8_0 , 
        \scalestate_0/fst_lst_pulse8_2 , 
        \scalestate_0/fst_lst_pulse8_9 , 
        \scalestate_0/fst_lst_pulse8_NE_4 , 
        \scalestate_0/necount[4]_net_1 , 
        \scalestate_0/NE_NUM[4]_net_1 , 
        \scalestate_0/fst_lst_pulse8_10 , 
        \scalestate_0/fst_lst_pulse8_NE_3 , 
        \scalestate_0/necount[8]_net_1 , 
        \scalestate_0/NE_NUM[8]_net_1 , 
        \scalestate_0/fst_lst_pulse8_7 , 
        \scalestate_0/necount[3]_net_1 , 
        \scalestate_0/NE_NUM[3]_net_1 , 
        \scalestate_0/fst_lst_pulse8_1 , 
        \scalestate_0/necount[6]_net_1 , 
        \scalestate_0/NE_NUM[6]_net_1 , 
        \scalestate_0/fst_lst_pulse8_5 , \scalestate_0/M_pulse8_NE_8 , 
        \scalestate_0/M_pulse8_NE_2 , \scalestate_0/M_pulse8_NE_1 , 
        \scalestate_0/M_pulse8_NE_5 , \scalestate_0/M_pulse8_0 , 
        \scalestate_0/M_pulse8_2 , \scalestate_0/M_pulse8_9 , 
        \scalestate_0/M_pulse8_NE_4 , \scalestate_0/M_NUM[4]_net_1 , 
        \scalestate_0/M_pulse8_10 , \scalestate_0/M_pulse8_NE_3 , 
        \scalestate_0/M_NUM[8]_net_1 , \scalestate_0/M_pulse8_7 , 
        \scalestate_0/M_NUM[3]_net_1 , \scalestate_0/M_pulse8_1 , 
        \scalestate_0/M_NUM[6]_net_1 , \scalestate_0/M_pulse8_5 , 
        \scalestate_0/un1_CS6_39_i_a3_1 , 
        \scalestate_0/un1_CS6_39_i_a3_0 , \scalestate_0/CS[6]_net_1 , 
        \scalestate_0/un1_CS6_17_i_a3_0 , \scalestate_0/CS[4]_net_1 , 
        \scalestate_0/un1_CS_44_i_0 , \scalestate_0/N_1212 , 
        \scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 , 
        \scalestate_0/un1_CS6_0 , \scalestate_0/CS[10]_net_1 , 
        \scalestate_0/CS[9]_net_1 , \scalestate_0/un1_CS6_39_i_a2_0 , 
        \scalestate_0/CS[18]_net_1 , \scalestate_0/un1_CS6_31_i_o2_0 , 
        \scalestate_0/CS[7]_net_1 , \scalestate_0/CS_RNO_1[2] , 
        \scalestate_0/un1_CS6_26 , \scalestate_0/M_pulse8_NE , 
        \scalestate_0/N_1304 , \scalestate_0/N_1097 , 
        \scalestate_0/N_1208 , \scalestate_0/timecount_20[21] , 
        \scalestate_0/OPENTIME_TEL_m[21] , 
        \scalestate_0/CS_RNO_0[8]_net_1 , \scalestate_0/un1_CS6 , 
        \scalestate_0/un1_CS6_34 , \scalestate_0/N_1309 , 
        \scalestate_0/sw_acq1_1_sqmuxa , \scalestate_0/N_258 , 
        \scalestate_0/fst_lst_pulse8_NE , \scalestate_0/un1_CS6_14 , 
        \scalestate_0/un1_CS_27 , \scalestate_0/intertodsp_1_sqmuxa , 
        \scalestate_0/N_1269 , \scalestate_0/N_1241 , 
        \scalestate_0/un1_CS_34 , \scalestate_0/N_1195 , 
        \scalestate_0/CS_i[0]_net_1 , 
        \scalestate_0/ACQ180_NUM_1_sqmuxa , \scalestate_0/N_67 , 
        \scalestate_0/N_62 , \scalestate_0/ACQ90_NUM_1_sqmuxa , 
        \scalestate_0/timecount_20[20] , 
        \scalestate_0/OPENTIME_TEL_m[20] , 
        \scalestate_0/timecount_16_sqmuxa_1 , \scalestate_0/N_543 , 
        \scalestate_0/N_1259 , \scalestate_0/N_544 , 
        \scalestate_0/N_723 , \scalestate_0/N_1167 , 
        \scalestate_0/N_727 , \scalestate_0/N_741 , 
        \scalestate_0/N_1181 , \scalestate_0/N_743 , 
        \scalestate_0/N_1163 , \scalestate_0/long_opentime_RNO_net_1 , 
        \scalestate_0/intertodsp_RNO_0_net_1 , 
        \scalestate_0/dump_start_RNO_0_net_1 , 
        \scalestate_0/rt_sw_RNO_1_net_1 , \scalestate_0/soft_d_RNO_2 , 
        \scalestate_0/necount_LE_NE_RNO_net_1 , 
        \scalestate_0/necount_LE_NE_1 , 
        \scalestate_0/necount_LE_M_RNO_net_1 , 
        \scalestate_0/necount_LE_M_1 , 
        \scalestate_0/fst_lst_pulse_RNO_net_1 , 
        \scalestate_0/strippluse_RNO[0]_net_1 , \scalestate_0/N_559 , 
        \scalestate_0/strippluse_RNO[1]_net_1 , \scalestate_0/N_560 , 
        \scalestate_0/strippluse_RNO[2]_net_1 , \scalestate_0/N_561 , 
        \scalestate_0/strippluse_RNO[3]_net_1 , \scalestate_0/N_562 , 
        \scalestate_0/strippluse_RNO[4]_net_1 , \scalestate_0/N_563 , 
        \scalestate_0/strippluse_RNO[5]_net_1 , \scalestate_0/N_564 , 
        \scalestate_0/strippluse_RNO[6]_net_1 , \scalestate_0/N_565 , 
        \scalestate_0/strippluse_RNO[7]_net_1 , \scalestate_0/N_566 , 
        \scalestate_0/strippluse_RNO[8]_net_1 , \scalestate_0/N_567 , 
        \scalestate_0/strippluse_RNO[9]_net_1 , \scalestate_0/N_568 , 
        \scalestate_0/strippluse_RNO[10]_net_1 , \scalestate_0/N_569 , 
        \scalestate_0/strippluse_RNO[11]_net_1 , \scalestate_0/N_570 , 
        \scalestate_0/s_acqnum_1_RNO[0]_net_1 , \scalestate_0/N_547 , 
        \scalestate_0/s_acqnum_1_RNO[1]_net_1 , \scalestate_0/N_548 , 
        \scalestate_0/s_acqnum_1_RNO[2]_net_1 , \scalestate_0/N_549 , 
        \scalestate_0/s_acqnum_1_RNO[3]_net_1 , \scalestate_0/N_550 , 
        \scalestate_0/s_acqnum_1_RNO[4]_net_1 , \scalestate_0/N_551 , 
        \scalestate_0/s_acqnum_1_RNO[5]_net_1 , \scalestate_0/N_552 , 
        \scalestate_0/s_acqnum_1_RNO[6]_net_1 , \scalestate_0/N_553 , 
        \scalestate_0/s_acqnum_1_RNO[7]_net_1 , \scalestate_0/N_554 , 
        \scalestate_0/s_acqnum_1_RNO[8]_net_1 , \scalestate_0/N_555 , 
        \scalestate_0/s_acqnum_1_RNO[9]_net_1 , \scalestate_0/N_556 , 
        \scalestate_0/s_acqnum_1_RNO[10]_net_1 , \scalestate_0/N_557 , 
        \scalestate_0/s_acqnum_1_RNO[11]_net_1 , \scalestate_0/N_558 , 
        \scalestate_0/s_acqnum_7[0] , \scalestate_0/s_acqnum_7[1] , 
        \scalestate_0/s_acqnum_7[2] , \scalestate_0/s_acqnum_7[3] , 
        \scalestate_0/s_acqnum_7[4] , \scalestate_0/s_acqnum_7[5] , 
        \scalestate_0/s_acqnum_7[6] , \scalestate_0/s_acqnum_7[7] , 
        \scalestate_0/s_acqnum_7[8] , \scalestate_0/s_acqnum_7[9] , 
        \scalestate_0/s_acqnum_7[10] , \scalestate_0/s_acqnum_7[11] , 
        \scalestate_0/strippluse_6[0] , \scalestate_0/strippluse_6[1] , 
        \scalestate_0/strippluse_6[2] , \scalestate_0/strippluse_6[3] , 
        \scalestate_0/strippluse_6[4] , \scalestate_0/strippluse_6[5] , 
        \scalestate_0/strippluse_6[6] , \scalestate_0/strippluse_6[7] , 
        \scalestate_0/strippluse_6[8] , \scalestate_0/strippluse_6[9] , 
        \scalestate_0/strippluse_6[10] , 
        \scalestate_0/strippluse_6[11] , 
        \scalestate_0/NE_NUM[0]_net_1 , 
        \scalestate_0/necount[0]_net_1 , 
        \scalestate_0/NE_NUM[1]_net_1 , 
        \scalestate_0/necount[1]_net_1 , 
        \scalestate_0/NE_NUM[2]_net_1 , 
        \scalestate_0/necount[2]_net_1 , 
        \scalestate_0/NE_NUM[5]_net_1 , 
        \scalestate_0/necount[5]_net_1 , 
        \scalestate_0/NE_NUM[7]_net_1 , 
        \scalestate_0/necount[7]_net_1 , 
        \scalestate_0/NE_NUM[9]_net_1 , 
        \scalestate_0/necount[9]_net_1 , 
        \scalestate_0/NE_NUM[10]_net_1 , 
        \scalestate_0/necount[10]_net_1 , \scalestate_0/N_431 , 
        \scalestate_0/STRIPNUM180_NUM[11]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[11]_net_1 , \scalestate_0/N_452 , 
        \scalestate_0/ACQ180_NUM[4]_net_1 , 
        \scalestate_0/ACQ90_NUM[4]_net_1 , \scalestate_0/N_453 , 
        \scalestate_0/ACQ180_NUM[5]_net_1 , 
        \scalestate_0/ACQ90_NUM[5]_net_1 , \scalestate_0/N_454 , 
        \scalestate_0/ACQ180_NUM[6]_net_1 , 
        \scalestate_0/ACQ90_NUM[6]_net_1 , \scalestate_0/N_455 , 
        \scalestate_0/ACQ180_NUM[7]_net_1 , 
        \scalestate_0/ACQ90_NUM[7]_net_1 , \scalestate_0/N_456 , 
        \scalestate_0/ACQ180_NUM[8]_net_1 , 
        \scalestate_0/ACQ90_NUM[8]_net_1 , 
        \scalestate_0/ACQECHO_NUM[4]_net_1 , 
        \scalestate_0/ACQECHO_NUM[5]_net_1 , 
        \scalestate_0/ACQECHO_NUM[6]_net_1 , 
        \scalestate_0/ACQECHO_NUM[7]_net_1 , 
        \scalestate_0/ACQECHO_NUM[8]_net_1 , 
        \scalestate_0/CS[11]_net_1 , \scalestate_0/N_1225 , 
        \scalestate_0/CS_RNO[14]_net_1 , \scalestate_0/N_1227 , 
        \scalestate_0/CS_RNO[16]_net_1 , \scalestate_0/N_1229 , 
        \scalestate_0/CS_RNO[20]_net_1 , \scalestate_0/N_1232 , 
        \scalestate_0/N_1203 , \scalestate_0/CS[17]_net_1 , 
        \scalestate_0/N_420 , \scalestate_0/STRIPNUM180_NUM[0]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[0]_net_1 , \scalestate_0/N_421 , 
        \scalestate_0/STRIPNUM180_NUM[1]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[1]_net_1 , \scalestate_0/N_422 , 
        \scalestate_0/STRIPNUM180_NUM[2]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[2]_net_1 , \scalestate_0/N_423 , 
        \scalestate_0/STRIPNUM180_NUM[3]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[3]_net_1 , \scalestate_0/N_424 , 
        \scalestate_0/STRIPNUM180_NUM[4]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[4]_net_1 , \scalestate_0/N_425 , 
        \scalestate_0/STRIPNUM180_NUM[5]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[5]_net_1 , \scalestate_0/N_426 , 
        \scalestate_0/STRIPNUM180_NUM[6]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[6]_net_1 , \scalestate_0/N_427 , 
        \scalestate_0/STRIPNUM180_NUM[7]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[7]_net_1 , \scalestate_0/N_428 , 
        \scalestate_0/STRIPNUM180_NUM[8]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[8]_net_1 , \scalestate_0/N_429 , 
        \scalestate_0/STRIPNUM180_NUM[9]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[9]_net_1 , \scalestate_0/N_430 , 
        \scalestate_0/STRIPNUM180_NUM[10]_net_1 , 
        \scalestate_0/STRIPNUM90_NUM[10]_net_1 , \scalestate_0/N_448 , 
        \scalestate_0/ACQ180_NUM[0]_net_1 , 
        \scalestate_0/ACQ90_NUM[0]_net_1 , \scalestate_0/N_449 , 
        \scalestate_0/ACQ180_NUM[1]_net_1 , 
        \scalestate_0/ACQ90_NUM[1]_net_1 , \scalestate_0/N_450 , 
        \scalestate_0/ACQ180_NUM[2]_net_1 , 
        \scalestate_0/ACQ90_NUM[2]_net_1 , \scalestate_0/N_451 , 
        \scalestate_0/ACQ180_NUM[3]_net_1 , 
        \scalestate_0/ACQ90_NUM[3]_net_1 , \scalestate_0/N_457 , 
        \scalestate_0/ACQ180_NUM[9]_net_1 , 
        \scalestate_0/ACQ90_NUM[9]_net_1 , \scalestate_0/N_458 , 
        \scalestate_0/ACQ180_NUM[10]_net_1 , 
        \scalestate_0/ACQ90_NUM[10]_net_1 , \scalestate_0/N_459 , 
        \scalestate_0/ACQ180_NUM[11]_net_1 , 
        \scalestate_0/ACQ90_NUM[11]_net_1 , 
        \scalestate_0/ACQECHO_NUM[0]_net_1 , 
        \scalestate_0/ACQECHO_NUM[1]_net_1 , 
        \scalestate_0/ACQECHO_NUM[2]_net_1 , 
        \scalestate_0/ACQECHO_NUM[3]_net_1 , 
        \scalestate_0/ACQECHO_NUM[9]_net_1 , 
        \scalestate_0/ACQECHO_NUM[10]_net_1 , 
        \scalestate_0/ACQECHO_NUM[11]_net_1 , 
        \scalestate_0/PLUSETIME90[0]_net_1 , 
        \scalestate_0/S_DUMPTIME[0]_net_1 , 
        \scalestate_0/CUTTIME90[0]_net_1 , 
        \scalestate_0/PLUSETIME180[0]_net_1 , 
        \scalestate_0/OPENTIME_TEL[0]_net_1 , 
        \scalestate_0/OPENTIME[0]_net_1 , 
        \scalestate_0/ACQTIME[0]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[0]_net_1 , 
        \scalestate_0/CUTTIME180[0]_net_1 , 
        \scalestate_0/PLUSETIME90[1]_net_1 , 
        \scalestate_0/S_DUMPTIME[1]_net_1 , 
        \scalestate_0/CUTTIME90[1]_net_1 , 
        \scalestate_0/PLUSETIME180[1]_net_1 , 
        \scalestate_0/OPENTIME_TEL[1]_net_1 , 
        \scalestate_0/OPENTIME[1]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[1]_net_1 , 
        \scalestate_0/CUTTIME180[1]_net_1 , 
        \scalestate_0/CUTTIMEI90[2]_net_1 , 
        \scalestate_0/PLUSETIME90[2]_net_1 , 
        \scalestate_0/PLUSETIME180[2]_net_1 , 
        \scalestate_0/OPENTIME_TEL[2]_net_1 , 
        \scalestate_0/OPENTIME[2]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[2]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[2]_net_1 , 
        \scalestate_0/CUTTIMEI90[4]_net_1 , 
        \scalestate_0/PLUSETIME90[4]_net_1 , 
        \scalestate_0/DUMPTIME[4]_net_1 , 
        \scalestate_0/S_DUMPTIME[4]_net_1 , 
        \scalestate_0/CUTTIME90[4]_net_1 , 
        \scalestate_0/PLUSETIME180[4]_net_1 , 
        \scalestate_0/OPENTIME_TEL[4]_net_1 , 
        \scalestate_0/OPENTIME[4]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[4]_net_1 , 
        \scalestate_0/CUTTIMEI90[5]_net_1 , 
        \scalestate_0/PLUSETIME90[5]_net_1 , 
        \scalestate_0/CUTTIME90[5]_net_1 , 
        \scalestate_0/PLUSETIME180[5]_net_1 , 
        \scalestate_0/OPENTIME_TEL[5]_net_1 , 
        \scalestate_0/OPENTIME[5]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[5]_net_1 , 
        \scalestate_0/PLUSETIME90[6]_net_1 , 
        \scalestate_0/CUTTIME90[6]_net_1 , 
        \scalestate_0/PLUSETIME180[6]_net_1 , 
        \scalestate_0/OPENTIME_TEL[6]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[6]_net_1 , 
        \scalestate_0/CUTTIME180[6]_net_1 , 
        \scalestate_0/PLUSETIME90[8]_net_1 , 
        \scalestate_0/DUMPTIME[8]_net_1 , 
        \scalestate_0/S_DUMPTIME[8]_net_1 , 
        \scalestate_0/CUTTIME90[8]_net_1 , 
        \scalestate_0/PLUSETIME180[8]_net_1 , 
        \scalestate_0/OPENTIME_TEL[8]_net_1 , 
        \scalestate_0/OPENTIME[8]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[8]_net_1 , 
        \scalestate_0/PLUSETIME90[10]_net_1 , 
        \scalestate_0/DUMPTIME[10]_net_1 , 
        \scalestate_0/S_DUMPTIME[10]_net_1 , 
        \scalestate_0/CUTTIME90[10]_net_1 , 
        \scalestate_0/PLUSETIME180[10]_net_1 , 
        \scalestate_0/OPENTIME_TEL[10]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[10]_net_1 , 
        \scalestate_0/CUTTIME180[10]_net_1 , 
        \scalestate_0/CUTTIMEI90[11]_net_1 , 
        \scalestate_0/PLUSETIME90[11]_net_1 , 
        \scalestate_0/DUMPTIME[11]_net_1 , 
        \scalestate_0/S_DUMPTIME[11]_net_1 , 
        \scalestate_0/CUTTIME90[11]_net_1 , 
        \scalestate_0/PLUSETIME180[11]_net_1 , 
        \scalestate_0/OPENTIME_TEL[11]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[11]_net_1 , 
        \scalestate_0/CUTTIME180[11]_net_1 , 
        \scalestate_0/PLUSETIME90[12]_net_1 , 
        \scalestate_0/S_DUMPTIME[12]_net_1 , 
        \scalestate_0/CUTTIME90[12]_net_1 , 
        \scalestate_0/PLUSETIME180[12]_net_1 , 
        \scalestate_0/OPENTIME_TEL[12]_net_1 , 
        \scalestate_0/OPENTIME[12]_net_1 , 
        \scalestate_0/ACQTIME[12]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[12]_net_1 , 
        \scalestate_0/CUTTIME180[12]_net_1 , 
        \scalestate_0/PLUSETIME90[13]_net_1 , 
        \scalestate_0/S_DUMPTIME[13]_net_1 , 
        \scalestate_0/CUTTIME90[13]_net_1 , 
        \scalestate_0/PLUSETIME180[13]_net_1 , 
        \scalestate_0/OPENTIME_TEL[13]_net_1 , 
        \scalestate_0/OPENTIME[13]_net_1 , 
        \scalestate_0/ACQTIME[13]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[13]_net_1 , 
        \scalestate_0/CUTTIME180[13]_net_1 , 
        \scalestate_0/PLUSETIME90[14]_net_1 , 
        \scalestate_0/S_DUMPTIME[14]_net_1 , 
        \scalestate_0/CUTTIME90[14]_net_1 , 
        \scalestate_0/PLUSETIME180[14]_net_1 , 
        \scalestate_0/OPENTIME_TEL[14]_net_1 , 
        \scalestate_0/OPENTIME[14]_net_1 , 
        \scalestate_0/ACQTIME[14]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[14]_net_1 , 
        \scalestate_0/CUTTIME180[14]_net_1 , 
        \scalestate_0/PLUSETIME90[15]_net_1 , 
        \scalestate_0/CUTTIME90[15]_net_1 , 
        \scalestate_0/PLUSETIME180[15]_net_1 , 
        \scalestate_0/OPENTIME_TEL[15]_net_1 , 
        \scalestate_0/OPENTIME[15]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[15]_net_1 , 
        \scalestate_0/CUTTIME180[15]_net_1 , 
        \scalestate_0/CUTTIME90[16]_net_1 , 
        \scalestate_0/OPENTIME_TEL[16]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[16]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[16]_net_1 , 
        \scalestate_0/CUTTIME180[16]_net_1 , 
        \scalestate_0/CUTTIME90[17]_net_1 , 
        \scalestate_0/OPENTIME_TEL[17]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[17]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[17]_net_1 , 
        \scalestate_0/CUTTIME180[17]_net_1 , 
        \scalestate_0/CUTTIME90[18]_net_1 , 
        \scalestate_0/OPENTIME_TEL[18]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[18]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[18]_net_1 , 
        \scalestate_0/CUTTIME180[18]_net_1 , 
        \scalestate_0/CUTTIME90[19]_net_1 , 
        \scalestate_0/OPENTIME_TEL[19]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[19]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[19]_net_1 , 
        \scalestate_0/CUTTIME180[19]_net_1 , 
        \scalestate_0/CUTTIME90[20]_net_1 , 
        \scalestate_0/OPENTIME_TEL[20]_net_1 , 
        \scalestate_0/CUTTIME180_Tini[20]_net_1 , 
        \scalestate_0/CS_RNO_1[1] , \scalestate_0/N_1217 , 
        \scalestate_0/CS_RNO_1[3] , \scalestate_0/N_1218 , 
        \scalestate_0/CS_RNO[10]_net_1 , \scalestate_0/N_1224 , 
        \scalestate_0/CS_RNO[13]_net_1 , \scalestate_0/N_1237 , 
        \scalestate_0/CS_RNO[15]_net_1 , \scalestate_0/N_1228 , 
        \scalestate_0/CS_RNO[17]_net_1 , \scalestate_0/N_1230 , 
        \scalestate_0/CS_RNO[18]_net_1 , \scalestate_0/N_1213 , 
        \scalestate_0/CS_RNO[19]_net_1 , \scalestate_0/N_1231 , 
        \scalestate_0/CS_i_RNO_0[0] , \scalestate_0/CS[1]_net_1 , 
        \scalestate_0/CS[3]_net_1 , \scalestate_0/N_66 , 
        \scalestate_0/N_65 , \scalestate_0/N_64 , \scalestate_0/N_61 , 
        \scalestate_0/S_DUMPTIME_1_sqmuxa , \scalestate_0/N_60 , 
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa , 
        \scalestate_0/NE_NUM_1_sqmuxa , \scalestate_0/N_1645 , 
        \scalestate_0/N_1661 , \scalestate_0/N_1665 , 
        \scalestate_0/N_1681 , \scalestate_0/N_1685 , 
        \scalestate_0/N_1701 , \scalestate_0/N_1707 , 
        \scalestate_0/N_1723 , \scalestate_0/N_1729 , 
        \scalestate_0/N_1745 , \scalestate_0/N_1751 , 
        \scalestate_0/N_1767 , \scalestate_0/N_1773 , 
        \scalestate_0/N_1789 , \scalestate_0/ACQECHO_NUM_1_sqmuxa , 
        \scalestate_0/ACQTIME_1_sqmuxa , \scalestate_0/M_NUM_1_sqmuxa , 
        \scalestate_0/CUTTIME180_Tini[9]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[9]_net_1 , 
        \scalestate_0/ACQTIME[9]_net_1 , 
        \scalestate_0/OPENTIME[9]_net_1 , 
        \scalestate_0/OPENTIME_TEL[9]_net_1 , 
        \scalestate_0/PLUSETIME180[9]_net_1 , 
        \scalestate_0/CUTTIME90[9]_net_1 , 
        \scalestate_0/PLUSETIME90[9]_net_1 , 
        \scalestate_0/CUTTIMEI90[9]_net_1 , 
        \scalestate_0/load_out_RNO_net_1 , \scalestate_0/N_572 , 
        \scalestate_0/N_1165 , \scalestate_0/N_1236 , 
        \scalestate_0/CS[21]_net_1 , \scalestate_0/N_1226 , 
        \scalestate_0/N_1177 , \scalestate_0/CS_RNO[21]_net_1 , 
        \scalestate_0/CS_RNO[12]_net_1 , \scalestate_0/N_1220 , 
        \scalestate_0/N_1219 , \scalestate_0/N_1175 , 
        \scalestate_0/N_1262 , \scalestate_0/N_1173 , 
        \scalestate_0/CS_RNO_1[5] , \scalestate_0/CS_RNO_1[4] , 
        \scalestate_0/N_297 , \scalestate_0/sw_acq2_RNO_1 , 
        \scalestate_0/N_541 , \scalestate_0/sw_acq1_RNO_0_net_1 , 
        \scalestate_0/N_542 , \scalestate_0/off_test_RNO_1_net_1 , 
        \scalestate_0/N_726 , \scalestate_0/dds_conf_RNO_0_net_1 , 
        \scalestate_0/N_728 , \scalestate_0/bb_ch_RNO_net_1 , 
        \scalestate_0/N_729 , \scalestate_0/N_744 , 
        \scalestate_0/N_1183 , 
        \scalestate_0/dump_sustain_ctrl_RNO_net_1 , 
        \scalestate_0/CS_RNO_1[6] , \scalestate_0/N_1221 , 
        \scalestate_0/CS_RNO_1[7] , \scalestate_0/N_1222 , 
        \scalestate_0/N_724 , \scalestate_0/N_1169 , 
        \scalestate_0/s_acq_RNO_net_1 , \scalestate_0/N_1189 , 
        \scalestate_0/N_1171 , 
        \scalestate_0/CUTTIME180_Tini[21]_net_1 , 
        \scalestate_0/OPENTIME_TEL[21]_net_1 , 
        \scalestate_0/CUTTIME90[21]_net_1 , \scalestate_0/N_1223 , 
        \scalestate_0/CS_RNO_0[9]_net_1 , 
        \scalestate_0/reset_out_RNO_net_1 , \scalestate_0/N_540 , 
        \scalestate_0/pluse_start_RNO_0_net_1 , \scalestate_0/N_725 , 
        \scalestate_0/s_acq180_RNO_net_1 , \scalestate_0/N_742 , 
        \scalestate_0/tetw_pluse_RNO_1 , \scalestate_0/N_1187 , 
        \scalestate_0/dumpoff_ctr_RNO_2 , \scalestate_0/pn_out_4 , 
        \scalestate_0/N_571 , \scalestate_0/N_1191 , 
        \scalestate_0/pn_out_RNO_net_1 , 
        \scalestate_0/PLUSETIME180_1_sqmuxa , 
        \scalestate_0/DUMPTIME_1_sqmuxa , 
        \scalestate_0/PLUSETIME90_0_sqmuxa , 
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa , 
        \scalestate_0/CUTTIME180_Tini[7]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[7]_net_1 , 
        \scalestate_0/OPENTIME[7]_net_1 , 
        \scalestate_0/OPENTIME_TEL[7]_net_1 , 
        \scalestate_0/PLUSETIME180[7]_net_1 , 
        \scalestate_0/CUTTIME90[7]_net_1 , 
        \scalestate_0/PLUSETIME90[7]_net_1 , \scalestate_0/N_1179 , 
        \scalestate_0/M_NUM[10]_net_1 , \scalestate_0/M_NUM[9]_net_1 , 
        \scalestate_0/M_NUM[7]_net_1 , \scalestate_0/M_NUM[5]_net_1 , 
        \scalestate_0/M_NUM[2]_net_1 , \scalestate_0/M_NUM[1]_net_1 , 
        \scalestate_0/M_NUM[0]_net_1 , \scalestate_0/N_740 , 
        \scalestate_0/necount1[10] , \scalestate_0/N_739 , 
        \scalestate_0/necount1[9] , \scalestate_0/N_738 , 
        \scalestate_0/necount1[8] , \scalestate_0/N_737 , 
        \scalestate_0/necount1[7] , \scalestate_0/N_736 , 
        \scalestate_0/necount1[6] , \scalestate_0/N_735 , 
        \scalestate_0/necount1[5] , \scalestate_0/N_734 , 
        \scalestate_0/necount1[4] , \scalestate_0/N_733 , 
        \scalestate_0/necount1[3] , \scalestate_0/N_732 , 
        \scalestate_0/necount1[2] , \scalestate_0/N_731 , 
        \scalestate_0/necount1[1] , 
        \scalestate_0/necount_RNO[0]_net_1 , 
        \scalestate_0/necount_RNO[10]_net_1 , 
        \scalestate_0/necount_RNO[9]_net_1 , 
        \scalestate_0/necount_RNO[8]_net_1 , 
        \scalestate_0/necount_RNO[7]_net_1 , 
        \scalestate_0/necount_RNO[6]_net_1 , 
        \scalestate_0/necount_RNO[5]_net_1 , 
        \scalestate_0/necount_RNO[4]_net_1 , 
        \scalestate_0/necount_RNO[3]_net_1 , 
        \scalestate_0/necount_RNO[2]_net_1 , 
        \scalestate_0/necount_RNO[1]_net_1 , 
        \scalestate_0/M_pulse_RNO_net_1 , \scalestate_0/N_745 , 
        \scalestate_0/CUTTIME180_Tini[3]_net_1 , 
        \scalestate_0/CUTTIME180_TEL[3]_net_1 , 
        \scalestate_0/OPENTIME[3]_net_1 , 
        \scalestate_0/OPENTIME_TEL[3]_net_1 , 
        \scalestate_0/PLUSETIME180[3]_net_1 , 
        \scalestate_0/PLUSETIME90[3]_net_1 , 
        \scalestate_0/CUTTIMEI90[3]_net_1 , 
        \scalestate_0/necount_cmp_0/OA1A_0_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_4_Y , 
        \scalestate_0/necount_cmp_0/NOR3A_2_Y , 
        \scalestate_0/necount_cmp_0/OR2A_4_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_5_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_6_Y , 
        \scalestate_0/necount_cmp_0/AND2A_0_Y , 
        \scalestate_0/necount_cmp_0/OR2A_1_Y , 
        \scalestate_0/necount_cmp_0/OA1C_0_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_7_Y , 
        \scalestate_0/necount_cmp_0/AO1_0_Y , 
        \scalestate_0/necount_cmp_0/AND2_0_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_1_Y , 
        \scalestate_0/necount_cmp_0/NOR3_0_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_0_Y , 
        \scalestate_0/necount_cmp_0/NOR3A_0_Y , 
        \scalestate_0/necount_cmp_0/OR2A_5_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_2_Y , 
        \scalestate_0/necount_cmp_0/OR2A_2_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_2_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_0_Y , 
        \scalestate_0/necount_cmp_0/OR2A_3_Y , 
        \scalestate_0/necount_cmp_0/AO1C_1_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_9_Y , 
        \scalestate_0/necount_cmp_0/AO1_1_Y , 
        \scalestate_0/necount_cmp_0/AND3_2_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_4_Y , 
        \scalestate_0/necount_cmp_0/NOR3A_1_Y , 
        \scalestate_0/necount_cmp_0/NAND3A_3_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_8_Y , 
        \scalestate_0/necount_cmp_0/AND3_1_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_5_Y , 
        \scalestate_0/necount_cmp_0/XNOR2_3_Y , 
        \scalestate_0/necount_cmp_0/OR2A_0_Y , 
        \scalestate_0/necount_cmp_0/AND3_0_Y , 
        \scalestate_0/necount_cmp_0/AO1C_0_Y , 
        \scalestate_0/necount_cmp_0/AO1C_2_Y , 
        \scalestate_0/necount_inc_0/Rcout_8_net , 
        \scalestate_0/necount_inc_0/Rcout_5_net , 
        \scalestate_0/necount_inc_0/inc_2_net , 
        \scalestate_0/necount_inc_0/inc_5_net , 
        \scalestate_0/necount_inc_0/Rcout_10_net , 
        \scalestate_0/necount_inc_0/inc_12_net , 
        \scalestate_0/necount_inc_0/inc_10_net , 
        \scalestate_0/necount_inc_0/Rcout_9_net , 
        \scalestate_0/necount_inc_0/incb_2_net , 
        \scalestate_0/necount_inc_0/inc_8_net , 
        \scalestate_0/necount_inc_0/Rcout_7_net , 
        \scalestate_0/necount_cmp_1/OA1A_0_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_4_Y , 
        \scalestate_0/necount_cmp_1/NOR3A_2_Y , 
        \scalestate_0/necount_cmp_1/OR2A_4_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_5_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_1_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_6_Y , 
        \scalestate_0/necount_cmp_1/AND2A_0_Y , 
        \scalestate_0/necount_cmp_1/OR2A_1_Y , 
        \scalestate_0/necount_cmp_1/OA1C_0_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_7_Y , 
        \scalestate_0/necount_cmp_1/AO1_0_Y , 
        \scalestate_0/necount_cmp_1/AND2_0_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_1_Y , 
        \scalestate_0/necount_cmp_1/NOR3_0_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_0_Y , 
        \scalestate_0/necount_cmp_1/NOR3A_0_Y , 
        \scalestate_0/necount_cmp_1/OR2A_5_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_2_Y , 
        \scalestate_0/necount_cmp_1/OR2A_2_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_0_Y , 
        \scalestate_0/necount_cmp_1/OR2A_3_Y , 
        \scalestate_0/necount_cmp_1/AO1C_1_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_9_Y , 
        \scalestate_0/necount_cmp_1/AO1_1_Y , 
        \scalestate_0/necount_cmp_1/AND3_2_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_4_Y , 
        \scalestate_0/necount_cmp_1/NOR3A_1_Y , 
        \scalestate_0/necount_cmp_1/NAND3A_3_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_8_Y , 
        \scalestate_0/necount_cmp_1/AND3_1_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_5_Y , 
        \scalestate_0/necount_cmp_1/XNOR2_3_Y , 
        \scalestate_0/necount_cmp_1/OR2A_0_Y , 
        \scalestate_0/necount_cmp_1/AND3_0_Y , 
        \scalestate_0/necount_cmp_1/AO1C_0_Y , 
        \scalestate_0/necount_cmp_1/AO1C_2_Y , 
        \topctrlchange_0/soft_dump_6 , \topctrlchange_0/s_dumpin2_m , 
        \topctrlchange_0/s_dumpin3_m , \topctrlchange_0/s_dumpin1_m , 
        \topctrlchange_0/un1_interin1[0] , 
        \topctrlchange_0/interin2_m , \topctrlchange_0/interin3_m , 
        \topctrlchange_0/interin1_m , \topctrlchange_0/N_8 , 
        \topctrlchange_0/N_10 , \topctrlchange_0/sw_acq1_6_iv , 
        \topctrlchange_0/N_12 , \topctrlchange_0/rt_sw_6 , 
        \topctrlchange_0/rt_sw_RNO_4 , 
        \topctrlchange_0/interupt_RNO_net_1 , 
        \topctrlchange_0/sw_acq1_RNO_1_net_1 , 
        \topctrlchange_0/rt_swin1_m , \topctrlchange_0/sw_acq1in3_i_m , 
        \topctrlchange_0/sw_acq2_6_iv , 
        \topctrlchange_0/sw_acq2in1_i_m , 
        \topctrlchange_0/sw_acq2_RNO_3 , \topctrlchange_0/N_9 , 
        \topctrlchange_0/soft_dump_RNO_0_net_1 , 
        \topctrlchange_0/N_11 , \GPMI_0/INV_0_Y , 
        \GPMI_0/xwe_xzcs2_syn_0/code_en_0_0 , 
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_net_1 , 
        \GPMI_0/xwe_xzcs2_syn_0/code_en_RNO_net_1 , 
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_net_1 , 
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_RNO_net_1 , 
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_RNO_net_1 , 
        \GPMI_0/rst_n_module_0/rst_nr2_net_1 , 
        \GPMI_0/rst_n_module_0/rst_nr1_net_1 , 
        \plusestate_0/CS_srsts_i_0[3] , \plusestate_0/CS[8]_net_1 , 
        \plusestate_0/CS_srsts_i_0[2] , \plusestate_0/CS[1]_net_1 , 
        \plusestate_0/CS_srsts_i_0[1] , \plusestate_0/CS_i[0]_net_1 , 
        \plusestate_0/CS_srsts_i_0[6] , \plusestate_0/CS[5]_net_1 , 
        \plusestate_0/CS_srsts_i_0[5] , \plusestate_0/CS[9]_net_1 , 
        \plusestate_0/CS_srsts_i_0[8] , \plusestate_0/CS[2]_net_1 , 
        \plusestate_0/CS_srsts_i_0[4] , \plusestate_0/CS[3]_net_1 , 
        \plusestate_0/CS_srsts_i_0[9] , \plusestate_0/CS[4]_net_1 , 
        \plusestate_0/timecount_cnst[3] , \plusestate_0/N_303 , 
        \plusestate_0/CS_RNO_0[1]_net_1 , 
        \plusestate_0/CS_RNO_0[2]_net_1 , 
        \plusestate_0/CS_RNO_0[3]_net_1 , 
        \plusestate_0/CS_RNO[8]_net_1 , 
        \plusestate_0/CS_RNO_0[4]_net_1 , 
        \plusestate_0/CS_RNO[9]_net_1 , 
        \plusestate_0/CS_RNO_0[5]_net_1 , \plusestate_0/N_298 , 
        \plusestate_0/N_302 , \plusestate_0/N_301 , 
        \plusestate_0/N_299 , \plusestate_0/CS_RNO_0[6]_net_1 , 
        \plusestate_0/CS[6]_net_1 , \plusestate_0/state_over_n_RNO_0 , 
        \plusestate_0/N_253 , \plusestate_0/N_247 , 
        \plusestate_0/N_245 , \plusestate_0/N_215 , 
        \plusestate_0/timecount_5[15] , \plusestate_0/N_86 , 
        \plusestate_0/N_271 , \plusestate_0/timecount_5[12] , 
        \plusestate_0/N_83 , \plusestate_0/timecount_5[10] , 
        \plusestate_0/N_81 , \plusestate_0/timecount_5[8] , 
        \plusestate_0/N_79 , \plusestate_0/timecount_5[7] , 
        \plusestate_0/N_78 , \plusestate_0/timecount_5[2] , 
        \plusestate_0/N_73 , \plusestate_0/timecount_5[1] , 
        \plusestate_0/N_72 , \plusestate_0/timecount_5[0] , 
        \plusestate_0/N_71 , \plusestate_0/DUMPTIME[15]_net_1 , 
        \plusestate_0/PLUSETIME[15]_net_1 , \plusestate_0/N_213 , 
        \plusestate_0/DUMPTIME[12]_net_1 , 
        \plusestate_0/PLUSETIME[12]_net_1 , 
        \plusestate_0/DUMPTIME[10]_net_1 , 
        \plusestate_0/PLUSETIME[10]_net_1 , 
        \plusestate_0/DUMPTIME[8]_net_1 , 
        \plusestate_0/PLUSETIME[8]_net_1 , 
        \plusestate_0/DUMPTIME[7]_net_1 , 
        \plusestate_0/PLUSETIME[7]_net_1 , 
        \plusestate_0/DUMPTIME[2]_net_1 , 
        \plusestate_0/PLUSETIME[2]_net_1 , 
        \plusestate_0/DUMPTIME[1]_net_1 , 
        \plusestate_0/PLUSETIME[1]_net_1 , 
        \plusestate_0/DUMPTIME[0]_net_1 , 
        \plusestate_0/PLUSETIME[0]_net_1 , \plusestate_0/CS_RNO_0[7] , 
        \plusestate_0/CS[7]_net_1 , 
        \plusestate_0/un1_sw_acq1_2_sqmuxa , 
        \plusestate_0/soft_d_RNO_1_net_1 , \plusestate_0/N_121 , 
        \plusestate_0/pluse_acq_RNO_net_1 , \plusestate_0/N_122 , 
        \plusestate_0/dds_config_RNO_net_1 , \plusestate_0/N_142 , 
        \plusestate_0/N_305 , \plusestate_0/N_141 , 
        \plusestate_0/off_test_RNO_0_net_1 , \plusestate_0/N_120 , 
        \plusestate_0/sw_acq1_RNO_net_1 , 
        \plusestate_0/DUMPTIME_1_sqmuxa_net_1 , 
        \plusestate_0/DUMPTIME_0_sqmuxa_net_1 , \plusestate_0/N_75 , 
        \plusestate_0/PLUSETIME[4]_net_1 , 
        \plusestate_0/DUMPTIME[4]_net_1 , \plusestate_0/N_76 , 
        \plusestate_0/PLUSETIME[5]_net_1 , 
        \plusestate_0/DUMPTIME[5]_net_1 , \plusestate_0/N_77 , 
        \plusestate_0/PLUSETIME[6]_net_1 , 
        \plusestate_0/DUMPTIME[6]_net_1 , \plusestate_0/N_80 , 
        \plusestate_0/PLUSETIME[9]_net_1 , 
        \plusestate_0/DUMPTIME[9]_net_1 , \plusestate_0/N_82 , 
        \plusestate_0/PLUSETIME[11]_net_1 , 
        \plusestate_0/DUMPTIME[11]_net_1 , \plusestate_0/N_84 , 
        \plusestate_0/PLUSETIME[13]_net_1 , 
        \plusestate_0/DUMPTIME[13]_net_1 , \plusestate_0/N_85 , 
        \plusestate_0/PLUSETIME[14]_net_1 , 
        \plusestate_0/DUMPTIME[14]_net_1 , 
        \plusestate_0/timecount_5[4] , \plusestate_0/N_249 , 
        \plusestate_0/timecount_5[5] , \plusestate_0/N_251 , 
        \plusestate_0/timecount_5[6] , \plusestate_0/N_223 , 
        \plusestate_0/timecount_5[9] , \plusestate_0/timecount_5[11] , 
        \plusestate_0/timecount_5[13] , \plusestate_0/timecount_5[14] , 
        \plusestate_0/tetw_pluse_RNO_0 , \plusestate_0/N_74 , 
        \plusestate_0/DUMPTIME[3]_net_1 , 
        \plusestate_0/PLUSETIME[3]_net_1 , 
        \plusestate_0/timecount_5[3] , 
        \plusestate_0/CS_i_RNO[0]_net_1 , 
        \bridge_div_0/clk_4f_reg1_net_1 , 
        \bridge_div_0/clk_4f_reg2_i_0 , 
        \bridge_div_0/count_RNIFNOM7[1]_net_1 , 
        \bridge_div_0/count_RNIEMOM7[0]_net_1 , 
        \bridge_div_0/count_RNIHPOM7[3]_net_1 , 
        \bridge_div_0/DWACT_FINC_E[0] , \bridge_div_0/clk_4f_reg1_i , 
        \bridge_div_0/un1_count_NE_1[0] , 
        \bridge_div_0/count[2]_net_1 , \bridge_div_0/dataall[2]_net_1 , 
        \bridge_div_0/un1_count_1_0[0] , 
        \bridge_div_0/un1_count_NE_0[0] , 
        \bridge_div_0/count[5]_net_1 , \bridge_div_0/count[4]_net_1 , 
        \bridge_div_0/un1_count_3[0] , 
        \bridge_div_0/clear1_n17_NE_1[0] , 
        \bridge_div_0/datahalf[2]_net_1 , 
        \bridge_div_0/clear1_n17_1[0] , 
        \bridge_div_0/clear1_n17_NE_0[0] , 
        \bridge_div_0/count[3]_net_1 , \bridge_div_0/un1_count_i[0] , 
        \bridge_div_0/un1_count_0[0] , \bridge_div_0/clear1_n17_NE[0] , 
        \bridge_div_0/clear1_n17_0[0] , \bridge_div_0/clk_4f_1_sqmuxa , 
        \bridge_div_0/dataall[3]_net_1 , 
        \bridge_div_0/datahalf[1]_net_1 , 
        \bridge_div_0/count[1]_net_1 , \bridge_div_0/dataall[1]_net_1 , 
        \bridge_div_0/datahalf[0]_net_1 , 
        \bridge_div_0/count[0]_net_1 , \bridge_div_0/dataall[0]_net_1 , 
        \bridge_div_0/count_RNIJROM7[5]_net_1 , 
        \bridge_div_0/clear1_n18 , 
        \bridge_div_0/count_RNIIQOM7[4]_net_1 , 
        \bridge_div_0/count_RNIGOOM7[2]_net_1 , 
        \bridge_div_0/clk_4f_5 , \bridge_div_0/clk_4f , 
        \bridge_div_0/DWACT_ADD_CI_0_partial_sum[0] , 
        \bridge_div_0/dataall_1[1] , \bridge_div_0/dataall_1[2] , 
        \bridge_div_0/dataall_1[3] , \bridge_div_0/count_5[0] , 
        \bridge_div_0/count_5[1] , \bridge_div_0/count_5[2] , 
        \bridge_div_0/count_5[3] , \bridge_div_0/count_5[4] , 
        \bridge_div_0/count_5[5] , \bridge_div_0/N_2 , 
        \bridge_div_0/N_4 , 
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0_1[0] , 
        \bridge_div_0/DWACT_ADD_CI_0_g_array_1[0] , 
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_2[0] , 
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0[0] , 
        \bridge_div_0/DWACT_ADD_CI_0_TMP[0] , 
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_1[0] , 
        \s_acq_change_0/s_load_0_0_RNIEJ0I1_net_1 , 
        \s_acq_change_0/s_rst_net_1 , \s_acq_change_0/s_stripnum_5[0] , 
        \s_acq_change_0/s_stripnum_5[1] , 
        \s_acq_change_0/s_stripnum_5[2] , 
        \s_acq_change_0/s_stripnum_5[3] , 
        \s_acq_change_0/s_stripnum_5[4] , 
        \s_acq_change_0/s_stripnum_5[5] , 
        \s_acq_change_0/s_stripnum_5[6] , 
        \s_acq_change_0/s_stripnum_5[7] , 
        \s_acq_change_0/s_stripnum_5[8] , 
        \s_acq_change_0/s_stripnum_5[9] , 
        \s_acq_change_0/s_stripnum_5[10] , 
        \s_acq_change_0/s_stripnum_5[11] , 
        \s_acq_change_0/s_acqnum_RNO[0]_net_1 , \s_acq_change_0/N_70 , 
        \s_acq_change_0/s_acqnum_RNO[1]_net_1 , \s_acq_change_0/N_71 , 
        \s_acq_change_0/s_acqnum_RNO[2]_net_1 , \s_acq_change_0/N_72 , 
        \s_acq_change_0/s_acqnum_RNO[3]_net_1 , \s_acq_change_0/N_73 , 
        \s_acq_change_0/s_acqnum_RNO[4]_net_1 , \s_acq_change_0/N_74 , 
        \s_acq_change_0/s_acqnum_RNO[5]_net_1 , \s_acq_change_0/N_75 , 
        \s_acq_change_0/s_acqnum_RNO[7]_net_1 , \s_acq_change_0/N_77 , 
        \s_acq_change_0/s_acqnum_RNO[8]_net_1 , \s_acq_change_0/N_78 , 
        \s_acq_change_0/s_acqnum_RNO[9]_net_1 , \s_acq_change_0/N_79 , 
        \s_acq_change_0/s_acqnum_RNO[11]_net_1 , \s_acq_change_0/N_81 , 
        \s_acq_change_0/s_acqnum_RNO[13]_net_1 , \s_acq_change_0/N_83 , 
        \s_acq_change_0/s_acqnum_RNO[14]_net_1 , \s_acq_change_0/N_84 , 
        \s_acq_change_0/s_acqnum_RNO[15]_net_1 , \s_acq_change_0/N_85 , 
        \s_acq_change_0/s_stripnum_RNO[0]_net_1 , 
        \s_acq_change_0/N_56 , 
        \s_acq_change_0/s_stripnum_RNO[1]_net_1 , 
        \s_acq_change_0/N_57 , 
        \s_acq_change_0/s_stripnum_RNO[2]_net_1 , 
        \s_acq_change_0/N_58 , 
        \s_acq_change_0/s_stripnum_RNO[3]_net_1 , 
        \s_acq_change_0/N_59 , 
        \s_acq_change_0/s_stripnum_RNO[4]_net_1 , 
        \s_acq_change_0/N_60 , 
        \s_acq_change_0/s_stripnum_RNO[5]_net_1 , 
        \s_acq_change_0/N_61 , 
        \s_acq_change_0/s_stripnum_RNO[6]_net_1 , 
        \s_acq_change_0/N_62 , 
        \s_acq_change_0/s_stripnum_RNO[7]_net_1 , 
        \s_acq_change_0/N_63 , 
        \s_acq_change_0/s_stripnum_RNO[8]_net_1 , 
        \s_acq_change_0/N_64 , 
        \s_acq_change_0/s_stripnum_RNO[9]_net_1 , 
        \s_acq_change_0/N_65 , 
        \s_acq_change_0/s_stripnum_RNO[10]_net_1 , 
        \s_acq_change_0/N_66 , 
        \s_acq_change_0/s_stripnum_RNO[11]_net_1 , 
        \s_acq_change_0/N_67 , \s_acq_change_0/s_acqnum_5[0] , 
        \s_acq_change_0/s_acqnum_5[1] , \s_acq_change_0/s_acqnum_5[2] , 
        \s_acq_change_0/s_acqnum_5[3] , \s_acq_change_0/s_acqnum_5[4] , 
        \s_acq_change_0/s_acqnum_5[5] , \s_acq_change_0/s_acqnum_5[7] , 
        \s_acq_change_0/s_acqnum_5[8] , \s_acq_change_0/s_acqnum_5[9] , 
        \s_acq_change_0/s_acqnum_5[11] , 
        \s_acq_change_0/s_acqnum_5[13] , 
        \s_acq_change_0/s_acqnum_5[14] , 
        \s_acq_change_0/s_acqnum_5[15] , \s_acq_change_0/N_69 , 
        \s_acq_change_0/s_load_5_net_1 , 
        \s_acq_change_0/s_rst_RNO_net_1 , \s_acq_change_0/N_68 , 
        \s_acq_change_0/s_rst_5 , \s_acq_change_0/s_acqnum_5[12] , 
        \s_acq_change_0/s_acqnum_5[10] , 
        \s_acq_change_0/s_acqnum_5[6] , \s_acq_change_0/N_82 , 
        \s_acq_change_0/N_80 , \s_acq_change_0/N_76 , 
        \s_acq_change_0/s_acqnum_RNO[12]_net_1 , 
        \s_acq_change_0/s_acqnum_RNO[10]_net_1 , 
        \s_acq_change_0/s_acqnum_RNO[6]_net_1 , \DUMP_0/count_2[0] , 
        \DUMP_0/count_2[1] , \DUMP_0/count_2[2] , \DUMP_0/count_2[3] , 
        \DUMP_0/count_2[4] , \DUMP_0/dump_state_0_off_start , 
        \DUMP_0/off_on_state_0_state_over , \DUMP_0/i[4] , 
        \DUMP_0/i[5] , \DUMP_0/i[6] , \DUMP_0/i[7] , \DUMP_0/i[8] , 
        \DUMP_0/i_2[0] , \DUMP_0/i_2[1] , \DUMP_0/i_0[2] , 
        \DUMP_0/i_0[3] , \DUMP_0/dump_state_0_timer_start , 
        \DUMP_0/dump_state_0_on_start , \DUMP_0/i_1[0] , 
        \DUMP_0/i_1[1] , \DUMP_0/i_0[0] , \DUMP_0/i_0[1] , 
        \DUMP_0/off_on_state_1_state_over , \DUMP_0/count[8] , 
        \DUMP_0/count[9] , \DUMP_0/count[10] , \DUMP_0/count[11] , 
        \DUMP_0/count_0[5] , \DUMP_0/count_0[6] , \DUMP_0/count_0[7] , 
        \DUMP_0/count_1[0] , \DUMP_0/count_1[1] , \DUMP_0/count_1[2] , 
        \DUMP_0/count_1[3] , \DUMP_0/count_1[4] , \DUMP_0/count_0[0] , 
        \DUMP_0/count_0[1] , \DUMP_0/count_0[2] , \DUMP_0/count_0[3] , 
        \DUMP_0/count_0[4] , 
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 , 
        \DUMP_0/off_on_timer_0/count_n4 , 
        \DUMP_0/off_on_timer_0/count_9_0 , 
        \DUMP_0/off_on_timer_0/count_n3 , 
        \DUMP_0/off_on_timer_0/count_c2 , 
        \DUMP_0/off_on_timer_0/count_n2 , 
        \DUMP_0/off_on_timer_0/count_c1 , 
        \DUMP_0/off_on_timer_0/count_n1 , 
        \DUMP_0/off_on_timer_0/count_n0 , 
        \DUMP_0/dump_state_0/un1_ns_0_a3_0 , 
        \DUMP_0/dump_state_0/N_206 , 
        \DUMP_0/dump_state_0/cs_RNO_1[5]_net_1 , 
        \DUMP_0/dump_state_0/N_1497_tz_tz , 
        \DUMP_0/dump_state_0/cs[6]_net_1 , \DUMP_0/dump_state_0/N_201 , 
        \DUMP_0/dump_state_0/cs_RNO_0[5]_net_1 , 
        \DUMP_0/dump_state_0/cs4 , \DUMP_0/dump_state_0/N_193 , 
        \DUMP_0/dump_state_0/N_167 , \DUMP_0/dump_state_0/N_203 , 
        \DUMP_0/dump_state_0/cs_RNO_0[4]_net_1 , 
        \DUMP_0/dump_state_0/N_185 , \DUMP_0/dump_state_0/N_186 , 
        \DUMP_0/dump_state_0/cs_RNO[2]_net_1 , 
        \DUMP_0/dump_state_0/N_182 , \DUMP_0/dump_state_0/N_183 , 
        \DUMP_0/dump_state_0/cs[4]_net_1 , 
        \DUMP_0/dump_state_0/cs_nsss[6] , \DUMP_0/dump_state_0/N_166 , 
        \DUMP_0/dump_state_0/N_176 , \DUMP_0/dump_state_0/N_196 , 
        \DUMP_0/dump_state_0/N_195 , \DUMP_0/dump_state_0/N_171 , 
        \DUMP_0/dump_state_0/N_173 , \DUMP_0/dump_state_0/ns[3] , 
        \DUMP_0/dump_state_0/cs[3]_net_1 , 
        \DUMP_0/dump_state_0/cs[1]_net_1 , 
        \DUMP_0/dump_state_0/cs_i_0[0]_net_1 , 
        \DUMP_0/dump_state_0/N_168 , \DUMP_0/dump_state_0/cs[7]_net_1 , 
        \DUMP_0/dump_state_0/off_start_RNO_net_1 , 
        \DUMP_0/dump_state_0/cs[2]_net_1 , 
        \DUMP_0/dump_state_0/cs_nsss[7] , 
        \DUMP_0/dump_state_0/cs_nsss[3] , 
        \DUMP_0/dump_state_0/cs_nsss[1] , 
        \DUMP_0/dump_state_0/timer_start_RNO_net_1 , 
        \DUMP_0/dump_state_0/N_88 , \DUMP_0/off_on_coder_1/i_0_2[1] , 
        \DUMP_0/off_on_coder_1/i_0_1[1] , 
        \DUMP_0/off_on_coder_1/i_RNO_1[1]_net_1 , 
        \DUMP_0/off_on_coder_1/i_RNO_1[0] , 
        \DUMP_0/off_on_state_1/N_36_i , \DUMP_0/off_on_state_1/N_42_i , 
        \DUMP_0/off_on_state_1/N_12_mux , \DUMP_0/off_on_state_1/N_10 , 
        \DUMP_0/off_on_state_1/cs[1]_net_1 , 
        \DUMP_0/off_on_state_1/N_9 , 
        \DUMP_0/off_on_state_1/cs_nsss[1] , 
        \DUMP_0/off_on_state_0/N_36_i , \DUMP_0/off_on_state_0/N_42_i , 
        \DUMP_0/off_on_state_0/N_12_mux , \DUMP_0/off_on_state_0/N_10 , 
        \DUMP_0/off_on_state_0/cs[1]_net_1 , 
        \DUMP_0/off_on_state_0/N_9 , 
        \DUMP_0/off_on_state_0/cs_nsss[1] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_12[3] , 
        \DUMP_0/dump_coder_0/un1_count_3_i[0] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_10[3] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE[0] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_7[3] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_6[3] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_8[3] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_5[3] , 
        \DUMP_0/dump_coder_0/un1_count_4_8[0] , 
        \DUMP_0/dump_coder_0/un1_count_4_9[0] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_3[3] , 
        \DUMP_0/dump_coder_0/un1_count_4_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_4_2[0] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_1[3] , 
        \DUMP_0/dump_coder_0/un1_count_4_10[0] , 
        \DUMP_0/dump_coder_0/un1_count_4_11[0] , 
        \DUMP_0/dump_coder_0/para1[7]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_4_6[0] , 
        \DUMP_0/dump_coder_0/para1[4]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_4_5[0] , 
        \DUMP_0/dump_coder_0/para1[0]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_4_1[0] , 
        \DUMP_0/dump_coder_0/i_0_0_a2_0[4] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_8[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_10[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_0_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_4[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_6[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_11[0] , 
        \DUMP_0/dump_coder_0/un1_count_2_NE_1[0] , 
        \DUMP_0/dump_coder_0/para3[9]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_2_8[0] , 
        \DUMP_0/dump_coder_0/para3[2]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_2_1[0] , 
        \DUMP_0/dump_coder_0/para3[6]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_2_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_8[0] , 
        \DUMP_0/dump_coder_0/un1_count_10[0] , 
        \DUMP_0/dump_coder_0/un1_count_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_4_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_6[0] , 
        \DUMP_0/dump_coder_0/un1_count_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_11[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE_1[0] , 
        \DUMP_0/dump_coder_0/para5[9]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_8[0] , 
        \DUMP_0/dump_coder_0/para5[2]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_1_0[0] , 
        \DUMP_0/dump_coder_0/para5[6]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_5[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_8[0] , 
        \DUMP_0/dump_coder_0/i_reg16_10[0] , 
        \DUMP_0/dump_coder_0/i_reg16_0[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_5[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_7[0] , 
        \DUMP_0/dump_coder_0/i_reg16_3[0] , 
        \DUMP_0/dump_coder_0/i_reg16_4[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_3[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_6[0] , 
        \DUMP_0/dump_coder_0/i_reg16_7[0] , 
        \DUMP_0/dump_coder_0/i_reg16_11[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE_1[0] , 
        \DUMP_0/dump_coder_0/para6[9]_net_1 , 
        \DUMP_0/dump_coder_0/i_reg16_8[0] , 
        \DUMP_0/dump_coder_0/para6[2]_net_1 , 
        \DUMP_0/dump_coder_0/i_reg16_1[0] , 
        \DUMP_0/dump_coder_0/para6[6]_net_1 , 
        \DUMP_0/dump_coder_0/i_reg16_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_8[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_10[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_0_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_4[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_6[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_11[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE_1[0] , 
        \DUMP_0/dump_coder_0/para4[9]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_1_8[0] , 
        \DUMP_0/dump_coder_0/para4[2]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_1_1[0] , 
        \DUMP_0/dump_coder_0/para4[6]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_1_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_8[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_10[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_0_0[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_5[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_4[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_3[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_6[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_7[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_11[0] , 
        \DUMP_0/dump_coder_0/un1_count_3_NE_1[0] , 
        \DUMP_0/dump_coder_0/para2[9]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_3_8[0] , 
        \DUMP_0/dump_coder_0/para2[2]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_3_1[0] , 
        \DUMP_0/dump_coder_0/para2[6]_net_1 , 
        \DUMP_0/dump_coder_0/un1_count_3_5[0] , 
        \DUMP_0/dump_coder_0/i_reg16_NE[0] , 
        \DUMP_0/dump_coder_0/un1_count_NE[0] , 
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] , 
        \DUMP_0/dump_coder_0/i_RNO[4]_net_1 , 
        \DUMP_0/dump_coder_0/N_19 , \DUMP_0/dump_coder_0/para15_net_1 , 
        \DUMP_0/dump_coder_0/para16_net_1 , 
        \DUMP_0/dump_coder_0/para17_net_1 , 
        \DUMP_0/dump_coder_0/para19_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO_0[3]_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO_0[1] , 
        \DUMP_0/dump_coder_0/i_RNO_0[2] , 
        \DUMP_0/dump_coder_0/para2[0]_net_1 , 
        \DUMP_0/dump_coder_0/para3[0]_net_1 , 
        \DUMP_0/dump_coder_0/para4[0]_net_1 , 
        \DUMP_0/dump_coder_0/para5[0]_net_1 , 
        \DUMP_0/dump_coder_0/para6[0]_net_1 , 
        \DUMP_0/dump_coder_0/para1[1]_net_1 , 
        \DUMP_0/dump_coder_0/para2[1]_net_1 , 
        \DUMP_0/dump_coder_0/para3[1]_net_1 , 
        \DUMP_0/dump_coder_0/para4[1]_net_1 , 
        \DUMP_0/dump_coder_0/para5[1]_net_1 , 
        \DUMP_0/dump_coder_0/para6[1]_net_1 , 
        \DUMP_0/dump_coder_0/para1[2]_net_1 , 
        \DUMP_0/dump_coder_0/para1[3]_net_1 , 
        \DUMP_0/dump_coder_0/para2[3]_net_1 , 
        \DUMP_0/dump_coder_0/para3[3]_net_1 , 
        \DUMP_0/dump_coder_0/para4[3]_net_1 , 
        \DUMP_0/dump_coder_0/para5[3]_net_1 , 
        \DUMP_0/dump_coder_0/para6[3]_net_1 , 
        \DUMP_0/dump_coder_0/para2[4]_net_1 , 
        \DUMP_0/dump_coder_0/para3[4]_net_1 , 
        \DUMP_0/dump_coder_0/para4[4]_net_1 , 
        \DUMP_0/dump_coder_0/para5[4]_net_1 , 
        \DUMP_0/dump_coder_0/para6[4]_net_1 , 
        \DUMP_0/dump_coder_0/para1[5]_net_1 , 
        \DUMP_0/dump_coder_0/para2[5]_net_1 , 
        \DUMP_0/dump_coder_0/para3[5]_net_1 , 
        \DUMP_0/dump_coder_0/para4[5]_net_1 , 
        \DUMP_0/dump_coder_0/para5[5]_net_1 , 
        \DUMP_0/dump_coder_0/para6[5]_net_1 , 
        \DUMP_0/dump_coder_0/para1[6]_net_1 , 
        \DUMP_0/dump_coder_0/para2[7]_net_1 , 
        \DUMP_0/dump_coder_0/para3[7]_net_1 , 
        \DUMP_0/dump_coder_0/para4[7]_net_1 , 
        \DUMP_0/dump_coder_0/para5[7]_net_1 , 
        \DUMP_0/dump_coder_0/para6[7]_net_1 , 
        \DUMP_0/dump_coder_0/para1[8]_net_1 , 
        \DUMP_0/dump_coder_0/para2[8]_net_1 , 
        \DUMP_0/dump_coder_0/para3[8]_net_1 , 
        \DUMP_0/dump_coder_0/para4[8]_net_1 , 
        \DUMP_0/dump_coder_0/para5[8]_net_1 , 
        \DUMP_0/dump_coder_0/para6[8]_net_1 , 
        \DUMP_0/dump_coder_0/para1[9]_net_1 , 
        \DUMP_0/dump_coder_0/para1[10]_net_1 , 
        \DUMP_0/dump_coder_0/para2[10]_net_1 , 
        \DUMP_0/dump_coder_0/para3[10]_net_1 , 
        \DUMP_0/dump_coder_0/para4[10]_net_1 , 
        \DUMP_0/dump_coder_0/para5[10]_net_1 , 
        \DUMP_0/dump_coder_0/para6[10]_net_1 , 
        \DUMP_0/dump_coder_0/para1[11]_net_1 , 
        \DUMP_0/dump_coder_0/para2[11]_net_1 , 
        \DUMP_0/dump_coder_0/para3[11]_net_1 , 
        \DUMP_0/dump_coder_0/para4[11]_net_1 , 
        \DUMP_0/dump_coder_0/para5[11]_net_1 , 
        \DUMP_0/dump_coder_0/para6[11]_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO[5]_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO[6]_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO[7]_net_1 , 
        \DUMP_0/dump_coder_0/i_RNO[8]_net_1 , 
        \DUMP_0/dump_coder_0/para18_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 , 
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 , 
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[0]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[1]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[2]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[3]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[4]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[5]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[6]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[7]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[8]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[9]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[10]_net_1 , 
        \DUMP_0/dump_coder_0/para2_4[11]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[0]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[1]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[2]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[3]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[4]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[5]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[6]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[7]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[8]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[9]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[10]_net_1 , 
        \DUMP_0/dump_coder_0/para4_4[11]_net_1 , 
        \DUMP_0/dump_coder_0/para5_4[0] , 
        \DUMP_0/dump_coder_0/para5_4[1] , 
        \DUMP_0/dump_coder_0/para5_4[2] , 
        \DUMP_0/dump_coder_0/para5_4[3] , 
        \DUMP_0/dump_coder_0/para5_4[4] , 
        \DUMP_0/dump_coder_0/para5_4[5] , 
        \DUMP_0/dump_coder_0/para5_4[6] , 
        \DUMP_0/dump_coder_0/para5_4[7] , 
        \DUMP_0/dump_coder_0/para5_4[8] , 
        \DUMP_0/dump_coder_0/para5_4[9] , 
        \DUMP_0/dump_coder_0/para5_4[10] , 
        \DUMP_0/dump_coder_0/para5_4[11] , 
        \DUMP_0/dump_coder_0/i_RNO_0[0] , \DUMP_0/dump_timer_0/N_52 , 
        \DUMP_0/dump_timer_0/count_c8 , 
        \DUMP_0/dump_timer_0/count_23_0 , 
        \DUMP_0/dump_timer_0/count_n10 , 
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 , 
        \DUMP_0/dump_timer_0/count_n10_tz , 
        \DUMP_0/dump_timer_0/count_c1 , \DUMP_0/dump_timer_0/count_c2 , 
        \DUMP_0/dump_timer_0/count_c3 , \DUMP_0/dump_timer_0/count_c4 , 
        \DUMP_0/dump_timer_0/count_c5 , \DUMP_0/dump_timer_0/count_c6 , 
        \DUMP_0/dump_timer_0/count_c7 , 
        \DUMP_0/dump_timer_0/count_n11 , 
        \DUMP_0/dump_timer_0/count_n2 , \DUMP_0/dump_timer_0/count_n3 , 
        \DUMP_0/dump_timer_0/count_n4 , \DUMP_0/dump_timer_0/count_n5 , 
        \DUMP_0/dump_timer_0/count_n6 , \DUMP_0/dump_timer_0/count_n7 , 
        \DUMP_0/dump_timer_0/count_n8 , \DUMP_0/dump_timer_0/count_n9 , 
        \DUMP_0/dump_timer_0/count_n0 , \DUMP_0/dump_timer_0/count_n1 , 
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 , 
        \DUMP_0/off_on_timer_1/count_n2 , 
        \DUMP_0/off_on_timer_1/count_c1 , 
        \DUMP_0/off_on_timer_1/count_n3 , 
        \DUMP_0/off_on_timer_1/count_c2 , 
        \DUMP_0/off_on_timer_1/count_n4 , 
        \DUMP_0/off_on_timer_1/count_9_0 , 
        \DUMP_0/off_on_timer_1/count_n0 , 
        \DUMP_0/off_on_timer_1/count_n1 , 
        \DUMP_0/off_on_coder_0/i_0_2[1] , 
        \DUMP_0/off_on_coder_0/i_0_1[1] , 
        \DUMP_0/off_on_coder_0/i_RNO_2[1] , 
        \DUMP_0/off_on_coder_0/i_RNO_2[0] , 
        \ClockManagement_0/clk_div500_0_clk_5K , 
        \ClockManagement_0/clk_5M_en , 
        \ClockManagement_0/pllclk_0_GLB , 
        \ClockManagement_0/long_timer_0/count_n11 , 
        \ClockManagement_0/long_timer_0/count_c10 , 
        \ClockManagement_0/long_timer_0/count[11]_net_1 , 
        \ClockManagement_0/long_timer_0/en_net_1 , 
        \ClockManagement_0/long_timer_0/count_c1 , 
        \ClockManagement_0/long_timer_0/count[1]_net_1 , 
        \ClockManagement_0/long_timer_0/count[0]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c2 , 
        \ClockManagement_0/long_timer_0/count[2]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c3 , 
        \ClockManagement_0/long_timer_0/count[3]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c4 , 
        \ClockManagement_0/long_timer_0/count[4]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c5 , 
        \ClockManagement_0/long_timer_0/count[5]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c6 , 
        \ClockManagement_0/long_timer_0/count[6]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c7 , 
        \ClockManagement_0/long_timer_0/count[7]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c8 , 
        \ClockManagement_0/long_timer_0/count[8]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c9 , 
        \ClockManagement_0/long_timer_0/count[10]_net_1 , 
        \ClockManagement_0/long_timer_0/count[9]_net_1 , 
        \ClockManagement_0/long_timer_0/count_m6_0_a2_7 , 
        \ClockManagement_0/long_timer_0/count_m6_0_a2_2 , 
        \ClockManagement_0/long_timer_0/count_m6_0_a2_1 , 
        \ClockManagement_0/long_timer_0/count_m6_0_a2_6 , 
        \ClockManagement_0/long_timer_0/count_m6_0_a2_4 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_13 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_2 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_1 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_10 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_12 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_0 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_7 , 
        \ClockManagement_0/long_timer_0/clear_n4_7 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_11 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_6 , 
        \ClockManagement_0/long_timer_0/clear_n4_8 , 
        \ClockManagement_0/long_timer_0/clear_n4_9 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_4 , 
        \ClockManagement_0/long_timer_0/clear_n4_1 , 
        \ClockManagement_0/long_timer_0/clear_n4_2 , 
        \ClockManagement_0/long_timer_0/clear_n4_5 , 
        \ClockManagement_0/long_timer_0/clear_n4_3 , 
        \ClockManagement_0/long_timer_0/clear_n4_6 , 
        \ClockManagement_0/long_timer_0/count[12]_net_1 , 
        \ClockManagement_0/long_timer_0/clear_n4_14 , 
        \ClockManagement_0/long_timer_0/clear_n4_13 , 
        \ClockManagement_0/long_timer_0/count[15]_net_1 , 
        \ClockManagement_0/long_timer_0/clk_5K_en_1 , 
        \ClockManagement_0/long_timer_0/count_c11 , 
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa , 
        \ClockManagement_0/long_timer_0/count_n15 , 
        \ClockManagement_0/long_timer_0/count_31_0 , 
        \ClockManagement_0/long_timer_0/count[14]_net_1 , 
        \ClockManagement_0/long_timer_0/count_c13 , 
        \ClockManagement_0/long_timer_0/count_n2 , 
        \ClockManagement_0/long_timer_0/count_n3 , 
        \ClockManagement_0/long_timer_0/count_n5 , 
        \ClockManagement_0/long_timer_0/count_n6 , 
        \ClockManagement_0/long_timer_0/count_n7 , 
        \ClockManagement_0/long_timer_0/count_n8 , 
        \ClockManagement_0/long_timer_0/count_n12 , 
        \ClockManagement_0/long_timer_0/count_n14 , 
        \ClockManagement_0/long_timer_0/count_n13 , 
        \ClockManagement_0/long_timer_0/count_c12 , 
        \ClockManagement_0/long_timer_0/count[13]_net_1 , 
        \ClockManagement_0/long_timer_0/count_n10 , 
        \ClockManagement_0/long_timer_0/count_n4 , 
        \ClockManagement_0/long_timer_0/count_n9 , 
        \ClockManagement_0/long_timer_0/N_95 , 
        \ClockManagement_0/long_timer_0/count_n1 , 
        \ClockManagement_0/long_timer_0/counte , 
        \ClockManagement_0/long_timer_0/timeup_RNO_net_1 , 
        \ClockManagement_0/long_timer_0/clk_5K_reg1_net_1 , 
        \ClockManagement_0/long_timer_0/clk_5K_reg2_net_1 , 
        \ClockManagement_0/long_timer_0/clk_5K_reg2_RNO_net_1 , 
        \ClockManagement_0/long_timer_0/clk_5K_reg1_RNO_net_1 , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_1[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_2[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_11[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_1_1[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_TMP[0] , 
        \ClockManagement_0/clk_div500_0/count[1]_net_1 , 
        \ClockManagement_0/clk_div500_0/count[6]_net_1 , 
        \ClockManagement_0/clk_div500_0/count[2]_net_1 , 
        \ClockManagement_0/clk_div500_0/count[4]_net_1 , 
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_6 , 
        \ClockManagement_0/clk_div500_0/count[0]_net_1 , 
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_5 , 
        \ClockManagement_0/clk_div500_0/count[5]_net_1 , 
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_2 , 
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_4 , 
        \ClockManagement_0/clk_div500_0/count[8]_net_1 , 
        \ClockManagement_0/clk_div500_0/count[3]_net_1 , 
        \ClockManagement_0/clk_div500_0/count[7]_net_1 , 
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa , 
        \ClockManagement_0/clk_div500_0/clk_5K_RNO_net_1 , 
        \ClockManagement_0/clk_div500_0/count_5[0] , 
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_partial_sum[0] , 
        \ClockManagement_0/clk_div500_0/count_5[8] , 
        \ClockManagement_0/clk_div500_0/I_38 , 
        \ClockManagement_0/clk_div500_0/count_5[7] , 
        \ClockManagement_0/clk_div500_0/I_36 , 
        \ClockManagement_0/clk_div500_0/count_5[6] , 
        \ClockManagement_0/clk_div500_0/I_34 , 
        \ClockManagement_0/clk_div500_0/count_5[5] , 
        \ClockManagement_0/clk_div500_0/I_32 , 
        \ClockManagement_0/clk_div500_0/count_5[4] , 
        \ClockManagement_0/clk_div500_0/I_31 , 
        \ClockManagement_0/clk_div500_0/count_5[3] , 
        \ClockManagement_0/clk_div500_0/I_37 , 
        \ClockManagement_0/clk_div500_0/count_5[2] , 
        \ClockManagement_0/clk_div500_0/I_35 , 
        \ClockManagement_0/clk_div500_0/count_5[1] , 
        \ClockManagement_0/clk_div500_0/I_33 , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_1[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_3[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_11[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_1[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_TMP[0] , 
        \ClockManagement_0/clk_10k_0/count[1]_net_1 , 
        \ClockManagement_0/clk_10k_0/count[6]_net_1 , 
        \ClockManagement_0/clk_10k_0/count[2]_net_1 , 
        \ClockManagement_0/clk_10k_0/count[4]_net_1 , 
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_6 , 
        \ClockManagement_0/clk_10k_0/count[7]_net_1 , 
        \ClockManagement_0/clk_10k_0/count[0]_net_1 , 
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_5 , 
        \ClockManagement_0/clk_10k_0/count[3]_net_1 , 
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_2 , 
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_4 , 
        \ClockManagement_0/clk_10k_0/count[8]_net_1 , 
        \ClockManagement_0/clk_10k_0/count[5]_net_1 , 
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa , 
        \ClockManagement_0/clk_10k_0/clk_5M_reg2_RNO_net_1 , 
        \ClockManagement_0/clk_10k_0/clk_5M_reg1_net_1 , 
        \ClockManagement_0/clk_10k_0/clk_5M_reg2_net_1 , 
        \ClockManagement_0/clk_10k_0/clk_5M_reg1_RNO_net_1 , 
        \ClockManagement_0/clk_10k_0/clock_10khz_RNO_net_1 , 
        \ClockManagement_0/clk_10k_0/clock_10khz_RNO_0_net_1 , 
        \ClockManagement_0/clk_10k_0/count_5[0] , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_partial_sum[0] , 
        \ClockManagement_0/clk_10k_0/count_5[8] , 
        \ClockManagement_0/clk_10k_0/I_38_0 , 
        \ClockManagement_0/clk_10k_0/count_5[7] , 
        \ClockManagement_0/clk_10k_0/I_36_0 , 
        \ClockManagement_0/clk_10k_0/count_5[6] , 
        \ClockManagement_0/clk_10k_0/I_34_0 , 
        \ClockManagement_0/clk_10k_0/count_5[5] , 
        \ClockManagement_0/clk_10k_0/I_32_0 , 
        \ClockManagement_0/clk_10k_0/count_5[4] , 
        \ClockManagement_0/clk_10k_0/I_31_0 , 
        \ClockManagement_0/clk_10k_0/count_5[3] , 
        \ClockManagement_0/clk_10k_0/I_37_0 , 
        \ClockManagement_0/clk_10k_0/count_5[2] , 
        \ClockManagement_0/clk_10k_0/I_35_0 , 
        \ClockManagement_0/clk_10k_0/count_5[1] , 
        \ClockManagement_0/clk_10k_0/I_33_0 , 
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_2[0] , 
        \DSTimer_0/AND2_0_Y , \DSTimer_0/net_0 , \DSTimer_0/DFI0_1_QN , 
        \DSTimer_0/dump_sustain_timer_0/start11_1 , 
        \DSTimer_0/dump_sustain_timer_0/count[2]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/data[2]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/un1_data_1 , 
        \DSTimer_0/dump_sustain_timer_0/start11_0 , 
        \DSTimer_0/dump_sustain_timer_0/count[3]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/data[3]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/enable_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/start11 , 
        \DSTimer_0/dump_sustain_timer_0/un1_data_0 , 
        \DSTimer_0/dump_sustain_timer_0/count_n2 , 
        \DSTimer_0/dump_sustain_timer_0/count_c1 , 
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p , 
        \DSTimer_0/dump_sustain_timer_0/count_n3 , 
        \DSTimer_0/dump_sustain_timer_0/count_7_0 , 
        \DSTimer_0/dump_sustain_timer_0/data_RNO[1]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/N_25 , 
        \DSTimer_0/dump_sustain_timer_0/data[1]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/data[0]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/count[1]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/count_n0 , 
        \DSTimer_0/dump_sustain_timer_0/count_n1 , 
        \DSTimer_0/dump_sustain_timer_0/N_27 , 
        \DSTimer_0/dump_sustain_timer_0/N_26 , 
        \DSTimer_0/dump_sustain_timer_0/N_24 , 
        \DSTimer_0/dump_sustain_timer_0/data_RNO[3]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/data_RNO[2]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/data_RNO[0]_net_1 , 
        \DSTimer_0/dump_sustain_timer_0/cmp_constant_4b_0/Temp_0_net , 
        \pd_pluse_top_0/i_0[4] , \pd_pluse_top_0/i_0[5] , 
        \pd_pluse_top_0/i_1[2] , \pd_pluse_top_0/i_1[3] , 
        \pd_pluse_top_0/i_6[0] , \pd_pluse_top_0/count[12] , 
        \pd_pluse_top_0/count[13] , \pd_pluse_top_0/count[14] , 
        \pd_pluse_top_0/count[15] , \pd_pluse_top_0/count_0[8] , 
        \pd_pluse_top_0/count_0[9] , \pd_pluse_top_0/count_0[10] , 
        \pd_pluse_top_0/count_0[11] , \pd_pluse_top_0/count_6[0] , 
        \pd_pluse_top_0/count_6[1] , \pd_pluse_top_0/count_6[2] , 
        \pd_pluse_top_0/count_6[3] , \pd_pluse_top_0/count_6[4] , 
        \pd_pluse_top_0/count_1[5] , \pd_pluse_top_0/count_1[6] , 
        \pd_pluse_top_0/count_1[7] , 
        \pd_pluse_top_0/pd_pluse_state_0_stateover , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_15[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_12[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_11[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_13[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_2[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_1[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_10[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_8[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_3[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_1[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_6[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_9[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_12[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_4[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_7[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_10[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[0]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_0[4] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[6]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_4[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[5]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_2[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[8]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_13[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[14]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_11[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[15]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_13[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_5[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_4[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_11[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_12[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_1[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_0[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_9[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_1[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_4[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_7[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_10[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_13[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_3[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[3]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_0[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[9]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_6[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[2]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_12[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[7]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_5[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[11]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_8[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[15]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_14[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_12[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_3[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_2[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_8[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_11[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_0[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_4[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_7[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_10[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_12[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_2[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_5[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_14[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_15[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_1[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[3]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_0[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[9]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_6[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[7]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_5[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[13]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_10[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[11]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_8[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_i[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa , 
        \pd_pluse_top_0/pd_pluse_coder_0/N_12 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[3] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[4]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_6[0] , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[0]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[0]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[1]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[1]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[1]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[2]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[2]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[3]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[4]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[4]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[4]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[5]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[5]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[6]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[6]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[7]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[8]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[8]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[9]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[10]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[10]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[10]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[11]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[12]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[12]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[12]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[13]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[13]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[14]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[14]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[15]_net_1 , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[2] , 
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[5] , 
        \pd_pluse_top_0/pd_pluse_state_0/en1_0_i_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_166 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_srsts_0_i_a5_1[12] , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[4]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[7]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[11]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[12]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_195 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[6]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_186 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_185 , 
        \pd_pluse_top_0/pd_pluse_state_0/en1_RNO_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_184 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[10]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_179 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_180 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[7]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/en2 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[3]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_174 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_175 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[8] , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_i[0]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[9]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_177 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_178 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[3]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[4] , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[11]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/stateover_RNO_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/en_RNO_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/en1_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[12]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_2[5] , 
        \pd_pluse_top_0/pd_pluse_state_0/N_187 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_176 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[2]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/N_173 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[1]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[5]_net_1 , 
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[1] , 
        \pd_pluse_top_0/pd_pluse_state_0/cs[8]_net_1 , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[0] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[1] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[1] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[2] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[2] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[3] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[3] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[4] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[4] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[5] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[5] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[6] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[6] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[7] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[7] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[8] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[8] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[9] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[9] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[10] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[10] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[11] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[11] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[12] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[12] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[13] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[13] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[14] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[14] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[15] , 
        \pd_pluse_top_0/pd_pluse_timer_0/count1[15] , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_8_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_5_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_13_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_20_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_14_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_10_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_12_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_11_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_14_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_9_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_22_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_5_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_15_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_8_net , 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_7_net , 
        \DUMP_ON_0/i_5[0] , \DUMP_ON_0/i_5[1] , 
        \DUMP_ON_0/off_on_state_0_state_over , \DUMP_ON_0/count_5[0] , 
        \DUMP_ON_0/count_5[1] , \DUMP_ON_0/count_5[2] , 
        \DUMP_ON_0/count_5[3] , \DUMP_ON_0/count_5[4] , 
        \DUMP_ON_0/off_on_state_0/N_36_i , 
        \DUMP_ON_0/off_on_state_0/N_42_i , 
        \DUMP_ON_0/off_on_state_0/cs_nsss[1] , 
        \DUMP_ON_0/off_on_state_0/N_10 , 
        \DUMP_ON_0/off_on_state_0/cs[1]_net_1 , 
        \DUMP_ON_0/off_on_state_0/N_9 , 
        \DUMP_ON_0/off_on_state_0/N_12_mux , 
        \DUMP_ON_0/off_on_coder_0/i_0_2[1] , 
        \DUMP_ON_0/off_on_coder_0/i_0_1[1] , 
        \DUMP_ON_0/off_on_coder_0/i_RNO_5[1] , 
        \DUMP_ON_0/off_on_coder_0/i_RNO_5[0] , 
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 , 
        \DUMP_ON_0/off_on_timer_0/count_n2 , 
        \DUMP_ON_0/off_on_timer_0/count_c1 , 
        \DUMP_ON_0/off_on_timer_0/count_n3 , 
        \DUMP_ON_0/off_on_timer_0/count_c2 , 
        \DUMP_ON_0/off_on_timer_0/count_n4 , 
        \DUMP_ON_0/off_on_timer_0/count_9_0 , 
        \DUMP_ON_0/off_on_timer_0/count_n0 , 
        \DUMP_ON_0/off_on_timer_0/count_n1 , 
        \nsctrl_choice_0/dumponoff_rst_5 , \nsctrl_choice_0/soft_d_5 , 
        \nsctrl_choice_0/soft_d_RNO_0_net_1 , 
        \nsctrl_choice_0/dumponoff_rst_RNO_net_1 , 
        \nsctrl_choice_0/dumpoff_ctr_RNO_1 , 
        \nsctrl_choice_0/dumpoff_ctr_5 , 
        \nsctrl_choice_0/sw_acq2_RNO_0_net_1 , 
        \nsctrl_choice_0/sw_acq2_5 , 
        \nsctrl_choice_0/intertodsp_RNO_net_1 , 
        \nsctrl_choice_0/intertodsp_5 , 
        \nsctrl_choice_0/rt_sw_RNO_0_net_1 , \nsctrl_choice_0/rt_sw_5 , 
        \nsctrl_choice_0/dumpon_ctr_5 , 
        \nsctrl_choice_0/dumpon_ctr_RNO_0_net_1 , 
        \scanstate_0/CS_srsts_i_0[1] , \scanstate_0/CS_li[0] , 
        \scanstate_0/CS_srsts_i_0[6] , \scanstate_0/CS[5]_net_1 , 
        \scanstate_0/CS_srsts_i_0[4] , \scanstate_0/CS[3]_net_1 , 
        \scanstate_0/CS_srsts_i_0[2] , \scanstate_0/CS[1]_net_1 , 
        \scanstate_0/CS_srsts_i_0[3] , \scanstate_0/CS[2]_net_1 , 
        \scanstate_0/CS_srsts_i_0[5] , \scanstate_0/CS[4]_net_1 , 
        \scanstate_0/CS_RNO_2[4] , \scanstate_0/CS_RNO_2[5] , 
        \scanstate_0/CS_RNO_2[3] , \scanstate_0/CS_RNO_2[2] , 
        \scanstate_0/timecount_cnst[4] , \scanstate_0/CS_RNO_2[1] , 
        \scanstate_0/CS_RNO_2[6] , \scanstate_0/CS[6]_net_1 , 
        \scanstate_0/N_111 , \scanstate_0/N_253 , 
        \scanstate_0/rt_sw_RNO_2 , 
        \scanstate_0/acqtime_0_sqmuxa_net_1 , 
        \scanstate_0/acqtime_1_sqmuxa_net_1 , \scanstate_0/N_59 , 
        \scanstate_0/acqtime[1]_net_1 , \scanstate_0/dectime[1]_net_1 , 
        \scanstate_0/N_194 , \scanstate_0/N_60 , 
        \scanstate_0/acqtime[2]_net_1 , \scanstate_0/dectime[2]_net_1 , 
        \scanstate_0/N_63 , \scanstate_0/acqtime[5]_net_1 , 
        \scanstate_0/dectime[5]_net_1 , \scanstate_0/N_64 , 
        \scanstate_0/acqtime[6]_net_1 , \scanstate_0/dectime[6]_net_1 , 
        \scanstate_0/N_65 , \scanstate_0/acqtime[7]_net_1 , 
        \scanstate_0/dectime[7]_net_1 , \scanstate_0/N_66 , 
        \scanstate_0/acqtime[8]_net_1 , \scanstate_0/dectime[8]_net_1 , 
        \scanstate_0/N_68 , \scanstate_0/acqtime[10]_net_1 , 
        \scanstate_0/dectime[10]_net_1 , \scanstate_0/N_70 , 
        \scanstate_0/acqtime[12]_net_1 , 
        \scanstate_0/dectime[12]_net_1 , \scanstate_0/N_71 , 
        \scanstate_0/acqtime[13]_net_1 , 
        \scanstate_0/dectime[13]_net_1 , \scanstate_0/N_72 , 
        \scanstate_0/acqtime[14]_net_1 , 
        \scanstate_0/dectime[14]_net_1 , \scanstate_0/timecount_5[2] , 
        \scanstate_0/timecount_cnst[2] , \scanstate_0/N_233 , 
        \scanstate_0/timecount_5[5] , \scanstate_0/timecount_5[6] , 
        \scanstate_0/timecount_5[7] , \scanstate_0/timecount_5[8] , 
        \scanstate_0/timecount_5[1] , \scanstate_0/timecount_5[10] , 
        \scanstate_0/timecount_5[12] , \scanstate_0/timecount_5[13] , 
        \scanstate_0/timecount_5[14] , \scanstate_0/CS_i_0_RNO_0[0] , 
        \scanstate_0/calctrl_RNO_net_1 , \scanstate_0/N_131 , 
        \scanstate_0/s_acq_RNO_0 , \scanstate_0/N_238 , 
        \scanstate_0/sw_acq2_RNO_2 , \scanstate_0/N_109 , 
        \scanstate_0/soft_d_RNO_3 , \scanstate_0/N_110 , 
        \scanstate_0/dds_conf_RNO_1 , \scanstate_0/N_130 , 
        \scanstate_0/CS_RNO_2[7] , \scanstate_0/CS[7]_net_1 , 
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa , 
        \scanstate_0/state_over_n_RNO_1 , \scanstate_0/N_255 , 
        \scanstate_0/dumpoff_ctr_RNO_3 , \scanstate_0/N_113 , 
        \scanstate_0/N_61 , \scanstate_0/dectime[3]_net_1 , 
        \scanstate_0/acqtime[3]_net_1 , \scanstate_0/N_67 , 
        \scanstate_0/dectime[9]_net_1 , \scanstate_0/acqtime[9]_net_1 , 
        \scanstate_0/N_69 , \scanstate_0/dectime[11]_net_1 , 
        \scanstate_0/acqtime[11]_net_1 , \scanstate_0/timecount_5[3] , 
        \scanstate_0/N_196 , \scanstate_0/timecount_5[9] , 
        \scanstate_0/timecount_5[11] , \scanstate_0/N_73 , 
        \scanstate_0/dectime[15]_net_1 , 
        \scanstate_0/acqtime[15]_net_1 , \scanstate_0/timecount_5[15] , 
        \scanstate_0/timecount_5[4] , \scanstate_0/N_62 , 
        \scanstate_0/timecount_5[0] , \scanstate_0/N_58 , 
        \scanstate_0/dectime[4]_net_1 , \scanstate_0/acqtime[4]_net_1 , 
        \scanstate_0/dectime[0]_net_1 , \scanstate_0/acqtime[0]_net_1 , 
        \DUMP_OFF_0/i_3[0] , \DUMP_OFF_0/i_3[1] , 
        \DUMP_OFF_0/off_on_state_0_state_over , 
        \DUMP_OFF_0/count_3[0] , \DUMP_OFF_0/count_3[1] , 
        \DUMP_OFF_0/count_3[2] , \DUMP_OFF_0/count_3[3] , 
        \DUMP_OFF_0/count_3[4] , \DUMP_OFF_0/off_on_state_0/N_36_i , 
        \DUMP_OFF_0/off_on_state_0/N_42_i , 
        \DUMP_OFF_0/off_on_state_0/N_12_mux , 
        \DUMP_OFF_0/off_on_state_0/N_10 , 
        \DUMP_OFF_0/off_on_state_0/cs[1]_net_1 , 
        \DUMP_OFF_0/off_on_state_0/N_9 , 
        \DUMP_OFF_0/off_on_state_0/cs_nsss[1] , 
        \DUMP_OFF_0/off_on_coder_0/i_0_2[1] , 
        \DUMP_OFF_0/off_on_coder_0/i_0_1[1] , 
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[1] , 
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[0] , 
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 , 
        \DUMP_OFF_0/off_on_timer_0/count_n2 , 
        \DUMP_OFF_0/off_on_timer_0/count_c1 , 
        \DUMP_OFF_0/off_on_timer_0/count_n3 , 
        \DUMP_OFF_0/off_on_timer_0/count_c2 , 
        \DUMP_OFF_0/off_on_timer_0/count_n4 , 
        \DUMP_OFF_0/off_on_timer_0/count_9_0 , 
        \DUMP_OFF_0/off_on_timer_0/count_n0 , 
        \DUMP_OFF_0/off_on_timer_0/count_n1 , 
        \n_acq_change_0/n_rst_n_0_net_1 , 
        \n_acq_change_0/n_acq_start_RNO_net_1 , 
        \n_acq_change_0/n_acq_start_5 , 
        \n_acq_change_0/n_rst_n_5_net_1 , 
        \noisestate_0/CS_srsts_i_0[6] , \noisestate_0/CS[5]_net_1 , 
        \noisestate_0/CS_srsts_i_0[5] , \noisestate_0/CS[4]_net_1 , 
        \noisestate_0/CS_srsts_i_0[2] , \noisestate_0/CS[1]_net_1 , 
        \noisestate_0/CS_srsts_i_0[3] , \noisestate_0/CS[2]_net_1 , 
        \noisestate_0/CS_srsts_i_0[4] , \noisestate_0/CS[3]_net_1 , 
        \noisestate_0/CS_srsts_i_0[1] , \noisestate_0/CS_li[0] , 
        \noisestate_0/CS_RNO[6]_net_1 , \noisestate_0/CS[6]_net_1 , 
        \noisestate_0/CS_RNO[5]_net_1 , \noisestate_0/CS_RNO[4]_net_1 , 
        \noisestate_0/CS_RNO[3]_net_1 , \noisestate_0/CS_RNO[1]_net_1 , 
        \noisestate_0/CS_RNO[2]_net_1 , 
        \noisestate_0/timecount_cnst[4] , 
        \noisestate_0/acqtime_0_sqmuxa_net_1 , 
        \noisestate_0/acqtime_1_sqmuxa_net_1 , \noisestate_0/N_57 , 
        \noisestate_0/acqtime[0]_net_1 , 
        \noisestate_0/dectime[0]_net_1 , \noisestate_0/N_191 , 
        \noisestate_0/N_58 , \noisestate_0/acqtime[1]_net_1 , 
        \noisestate_0/dectime[1]_net_1 , \noisestate_0/N_59 , 
        \noisestate_0/acqtime[2]_net_1 , 
        \noisestate_0/dectime[2]_net_1 , \noisestate_0/N_61 , 
        \noisestate_0/acqtime[4]_net_1 , 
        \noisestate_0/dectime[4]_net_1 , \noisestate_0/N_62 , 
        \noisestate_0/acqtime[5]_net_1 , 
        \noisestate_0/dectime[5]_net_1 , \noisestate_0/N_63 , 
        \noisestate_0/acqtime[6]_net_1 , 
        \noisestate_0/dectime[6]_net_1 , \noisestate_0/N_64 , 
        \noisestate_0/acqtime[7]_net_1 , 
        \noisestate_0/dectime[7]_net_1 , \noisestate_0/N_65 , 
        \noisestate_0/acqtime[8]_net_1 , 
        \noisestate_0/dectime[8]_net_1 , \noisestate_0/N_67 , 
        \noisestate_0/acqtime[10]_net_1 , 
        \noisestate_0/dectime[10]_net_1 , \noisestate_0/N_69 , 
        \noisestate_0/acqtime[12]_net_1 , 
        \noisestate_0/dectime[12]_net_1 , \noisestate_0/N_70 , 
        \noisestate_0/acqtime[13]_net_1 , 
        \noisestate_0/dectime[13]_net_1 , \noisestate_0/N_71 , 
        \noisestate_0/acqtime[14]_net_1 , 
        \noisestate_0/dectime[14]_net_1 , \noisestate_0/N_72 , 
        \noisestate_0/acqtime[15]_net_1 , 
        \noisestate_0/dectime[15]_net_1 , 
        \noisestate_0/timecount_5[0] , \noisestate_0/N_228 , 
        \noisestate_0/timecount_5[2] , 
        \noisestate_0/timecount_cnst[2] , 
        \noisestate_0/timecount_5[4] , \noisestate_0/timecount_5[5] , 
        \noisestate_0/timecount_5[6] , \noisestate_0/timecount_5[7] , 
        \noisestate_0/timecount_5[8] , \noisestate_0/timecount_5[1] , 
        \noisestate_0/timecount_5[10] , \noisestate_0/timecount_5[12] , 
        \noisestate_0/timecount_5[13] , \noisestate_0/timecount_5[14] , 
        \noisestate_0/timecount_5[15] , \noisestate_0/N_229 , 
        \noisestate_0/n_acq_RNO_net_1 , \noisestate_0/N_129 , 
        \noisestate_0/N_193 , \noisestate_0/timecount_5[11] , 
        \noisestate_0/N_68 , \noisestate_0/timecount_5[9] , 
        \noisestate_0/N_66 , \noisestate_0/timecount_5[3] , 
        \noisestate_0/N_60 , \noisestate_0/acqtime[11]_net_1 , 
        \noisestate_0/dectime[11]_net_1 , 
        \noisestate_0/acqtime[9]_net_1 , 
        \noisestate_0/dectime[9]_net_1 , 
        \noisestate_0/acqtime[3]_net_1 , 
        \noisestate_0/dectime[3]_net_1 , 
        \noisestate_0/soft_d_RNO_net_1 , \noisestate_0/N_109 , 
        \noisestate_0/dumpon_ctr_RNO_net_1 , \noisestate_0/N_130 , 
        \noisestate_0/N_248 , \noisestate_0/CS_RNO[7]_net_1 , 
        \noisestate_0/CS[7]_net_1 , 
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa , 
        \noisestate_0/state_over_n_RNO_net_1 , \noisestate_0/N_250 , 
        \noisestate_0/CS_i_0_RNO[0]_net_1 , \noisestate_0/N_233 , 
        \noisestate_0/sw_acq2_RNO_net_1 , \noisestate_0/N_108 , 
        \noisestate_0/rt_sw_RNO_net_1 , \noisestate_0/N_110 , 
        \noisestate_0/dumpoff_ctr_RNO_0_net_1 , \noisestate_0/N_112 , 
        \dds_change_0/dds_conf_6 , \dds_change_0/dds_confin2_m , 
        \dds_change_0/dds_confin3_m , \dds_change_0/dds_confin1_m , 
        \dds_change_0/dds_rst_6 , \dds_change_0/ddsrstin2_m , 
        \dds_change_0/ddsrstin3_m , \dds_change_0/ddsrstin1_m , 
        \dds_change_0/N_5 , \dds_change_0/N_6 , 
        \dds_change_0/dds_conf_RNO_net_1 , 
        \dds_change_0/dds_rst_RNO_net_1 , \xd_pad[6]/U0/NET1 , 
        \xd_pad[6]/U0/NET2 , \xd_pad[6]/U0/NET3 , \xa_pad[6]/U0/NET1 , 
        \soft_dump_pad/U0/NET1 , \soft_dump_pad/U0/NET2 , 
        \xa_pad[0]/U0/NET1 , \xd_pad[13]/U0/NET1 , 
        \xd_pad[13]/U0/NET2 , \xd_pad[13]/U0/NET3 , 
        \relay_on_pad[1]/U0/NET1 , \relay_on_pad[1]/U0/NET2 , 
        \xa_pad[5]/U0/NET1 , \ADC_pad[0]/U0/NET1 , 
        \xa_pad[12]/U0/NET1 , \relay_on_pad[0]/U0/NET1 , 
        \relay_on_pad[0]/U0/NET2 , \s_acq180_pad/U0/NET1 , 
        \s_acq180_pad/U0/NET2 , \relay_on_pad[5]/U0/NET1 , 
        \relay_on_pad[5]/U0/NET2 , \ddsfqud_pad/U0/NET1 , 
        \ddsfqud_pad/U0/NET2 , \gpio_pad/U0/NET1 , \Q2Q7_pad/U0/NET1 , 
        \Q2Q7_pad/U0/NET2 , \xd_pad[0]/U0/NET1 , \xd_pad[0]/U0/NET2 , 
        \xd_pad[0]/U0/NET3 , \ADC_pad[1]/U0/NET1 , 
        \ADC_pad[8]/U0/NET1 , \pulse_start_pad/U0/NET1 , 
        \pulse_start_pad/U0/NET2 , \xd_pad[9]/U0/NET1 , 
        \xd_pad[9]/U0/NET2 , \xd_pad[9]/U0/NET3 , 
        \interupt_pad/U0/NET1 , \interupt_pad/U0/NET2 , 
        \relay_close_pad[8]/U0/NET1 , \relay_close_pad[8]/U0/NET2 , 
        \sw_acq1_pad/U0/NET1 , \sw_acq1_pad/U0/NET2 , 
        \ADC_pad[9]/U0/NET1 , \Acq_clk_pad/U0/NET1 , 
        \Acq_clk_pad/U0/NET2 , \ADC_pad[2]/U0/NET1 , 
        \relay_close_pad[2]/U0/NET1 , \relay_close_pad[2]/U0/NET2 , 
        OCX40MHz_c, \dumpon_pad/U0/NET1 , \dumpon_pad/U0/NET2 , 
        \xa_pad[3]/U0/NET1 , \relay_on_pad[9]/U0/NET1 , 
        \relay_on_pad[9]/U0/NET2 , \k1_pad/U0/NET1 , \k1_pad/U0/NET2 , 
        \ddsreset_pad/U0/NET1 , \ddsreset_pad/U0/NET2 , 
        \sd_acq_en_pad/U0/NET1 , \sd_acq_en_pad/U0/NET2 , 
        \ADC_pad[11]/U0/NET1 , \xwe_pad/U0/NET1 , \xa_pad[10]/U0/NET1 , 
        \xd_pad[15]/U0/NET1 , \xd_pad[15]/U0/NET2 , 
        \xd_pad[15]/U0/NET3 , \ADC_pad[10]/U0/NET1 , 
        \xd_pad[7]/U0/NET1 , \xd_pad[7]/U0/NET2 , \xd_pad[7]/U0/NET3 , 
        \ddsdata_pad/U0/NET1 , \ddsdata_pad/U0/NET2 , 
        \xa_pad[11]/U0/NET1 , \Q1Q8_pad/U0/NET1 , \Q1Q8_pad/U0/NET2 , 
        \relay_on_pad[8]/U0/NET1 , \relay_on_pad[8]/U0/NET2 , 
        \dumpoff_pad/U0/NET1 , \dumpoff_pad/U0/NET2 , 
        \xa_pad[8]/U0/NET1 , \syn_md_out_pad/U0/NET1 , 
        \syn_md_out_pad/U0/NET2 , \ADC_pad[4]/U0/NET1 , 
        \relay_close_pad[9]/U0/NET1 , \relay_close_pad[9]/U0/NET2 , 
        \ADC_pad[3]/U0/NET1 , \XRD_pad/U0/NET1 , \xa_pad[4]/U0/NET1 , 
        \calcuinter_pad/U0/NET1 , \calcuinter_pad/U0/NET2 , 
        \relay_on_pad[7]/U0/NET1 , \relay_on_pad[7]/U0/NET2 , 
        \xa_pad[14]/U0/NET1 , \xd_pad[12]/U0/NET1 , 
        \xd_pad[12]/U0/NET2 , \xd_pad[12]/U0/NET3 , 
        \ddsclkout_pad/U0/NET1 , \relay_close_pad[0]/U0/NET1 , 
        \relay_close_pad[0]/U0/NET2 , \xa_pad[1]/U0/NET1 , 
        \xa_pad[2]/U0/NET1 , \relay_close_pad[7]/U0/NET1 , 
        \relay_close_pad[7]/U0/NET2 , \xa_pad[13]/U0/NET1 , 
        \xa_pad[7]/U0/NET1 , \xa_pad[17]/U0/NET1 , \GLA_pad/U0/NET1 , 
        \GLA_pad/U0/NET2 , \relay_close_pad[6]/U0/NET1 , 
        \relay_close_pad[6]/U0/NET2 , \xa_pad[16]/U0/NET1 , 
        \xa_pad[9]/U0/NET1 , \relay_on_pad[6]/U0/NET1 , 
        \relay_on_pad[6]/U0/NET2 , \rt_sw_pad/U0/NET1 , 
        \rt_sw_pad/U0/NET2 , \tri_ctrl_pad/U0/NET1 , 
        \relay_on_pad[3]/U0/NET1 , \relay_on_pad[3]/U0/NET2 , 
        \relay_close_pad[1]/U0/NET1 , \relay_close_pad[1]/U0/NET2 , 
        \k2_pad/U0/NET1 , \k2_pad/U0/NET2 , \sigtimeup_pad/U0/NET1 , 
        \sigtimeup_pad/U0/NET2 , \xd_pad[10]/U0/NET1 , 
        \xd_pad[10]/U0/NET2 , \xd_pad[10]/U0/NET3 , 
        \xa_pad[18]/U0/NET1 , \xd_pad[4]/U0/NET1 , \xd_pad[4]/U0/NET2 , 
        \xd_pad[4]/U0/NET3 , \ADC_pad[6]/U0/NET1 , 
        \pd_pulse_en_pad/U0/NET1 , \pd_pulse_en_pad/U0/NET2 , 
        \xd_pad[8]/U0/NET1 , \xd_pad[8]/U0/NET2 , \xd_pad[8]/U0/NET3 , 
        \relay_on_pad[2]/U0/NET1 , \relay_on_pad[2]/U0/NET2 , 
        \syn_md_tmp_pad/U0/NET1 , \syn_md_tmp_pad/U0/NET2 , 
        \xd_pad[1]/U0/NET1 , \xd_pad[1]/U0/NET2 , \xd_pad[1]/U0/NET3 , 
        \xd_pad[11]/U0/NET1 , \xd_pad[11]/U0/NET2 , 
        \xd_pad[11]/U0/NET3 , \zcs2_pad/U0/NET1 , \xd_pad[3]/U0/NET1 , 
        \xd_pad[3]/U0/NET2 , \xd_pad[3]/U0/NET3 , \ADC_pad[7]/U0/NET1 , 
        \ddswclk_pad/U0/NET1 , \ddswclk_pad/U0/NET2 , 
        \xa_pad[15]/U0/NET1 , \relay_on_pad[4]/U0/NET1 , 
        \relay_on_pad[4]/U0/NET2 , \relay_close_pad[5]/U0/NET1 , 
        \relay_close_pad[5]/U0/NET2 , \Q4Q5_pad/U0/NET1 , 
        \Q4Q5_pad/U0/NET2 , \xd_pad[5]/U0/NET1 , \xd_pad[5]/U0/NET2 , 
        \xd_pad[5]/U0/NET3 , \xd_pad[14]/U0/NET1 , 
        \xd_pad[14]/U0/NET2 , \xd_pad[14]/U0/NET3 , 
        \xd_pad[2]/U0/NET1 , \xd_pad[2]/U0/NET2 , \xd_pad[2]/U0/NET3 , 
        \relay_close_pad[4]/U0/NET1 , \relay_close_pad[4]/U0/NET2 , 
        \Q3Q6_pad/U0/NET1 , \Q3Q6_pad/U0/NET2 , \cal_out_pad/U0/NET1 , 
        \cal_out_pad/U0/NET2 , \relay_close_pad[3]/U0/NET1 , 
        \relay_close_pad[3]/U0/NET2 , \ADC_pad[5]/U0/NET1 , 
        \sw_acq2_pad/U0/NET1 , \sw_acq2_pad/U0/NET2 , 
        \PLUSE_0/bri_timer_0/count[5]/Y , 
        \PLUSE_0/bri_timer_0/count[6]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5]/Y , 
        \PLUSE_0/bri_timer_0/count[2]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10]/Y , 
        \PLUSE_0/bri_timer_0/count[4]/Y , \PLUSE_0/bri_coder_0/i[4]/Y , 
        \PLUSE_0/bri_coder_0/i[1]/Y , \PLUSE_0/bri_timer_0/count[7]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11]/Y , 
        \PLUSE_0/bri_coder_0/i[3]/Y , \PLUSE_0/bri_timer_0/count[1]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2]/Y , 
        \PLUSE_0/bri_coder_0/i[0]/Y , \PLUSE_0/bri_state_0/up/Y , 
        \bridge_div_0/clk_4f/Y , \PLUSE_0/bri_timer_0/count[3]/Y , 
        \PLUSE_0/bri_coder_0/i[2]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9]/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7]/Y , 
        \PLUSE_0/bri_state_0/down/Y , 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6]/Y , 
        AFLSDF_VCC, AFLSDF_GND;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[11]_net_1 ));
    MX2 \scalestate_0/strippluse_RNO_0[2]  (.A(
        \scalestate_0/strippluse_6[2] ), .B(
        \scalestate_0_strippluse[2] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_561 ));
    NOR2A \DUMP_0/dump_timer_0/count_RNO[0]  (.A(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_0/count_1[0] ), .Y(\DUMP_0/dump_timer_0/count_n0 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[26]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[26]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_470 ));
    DFN1E1 \state_1ms_0/PLUSETIME[5]  (.D(
        \top_code_0_state_1ms_data[5] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[5]_net_1 ));
    OA1C \top_code_0/n_rd_en_RNO  (.A(\top_code_0/N_207 ), .B(
        top_code_0_n_rd_en), .C(\top_code_0/N_282 ), .Y(
        \top_code_0/N_74 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[13]_net_1 )
        );
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_2  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] )
        );
    NOR2B \state_1ms_0/timecount_RNO_6[8]  (.A(
        \state_1ms_0/PLUSETIME[8]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[8] ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNIO1MJ[7]  (.A(
        \DUMP_0/dump_coder_0/para5[7]_net_1 ), .B(\DUMP_0/count_0[7] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_7[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[28]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[28]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_479 ));
    DFN1 \PLUSE_0/qq_timer_0/count[4]  (.D(
        \PLUSE_0/qq_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_9[4] ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[15]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO[15]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/sd_sacq_state_0/cs[15]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO[4]  (.A(\noisestate_0/N_61 ), .B(
        \noisestate_0/timecount_cnst[4] ), .S(\noisestate_0/N_228 ), 
        .Y(\noisestate_0/timecount_5[4] ));
    NOR3B \scalestate_0/timecount_ret_33_RNO  (.A(
        \scalestate_0/timecount_m1_e_2_0 ), .B(\scalestate_0/N_1089 ), 
        .C(\scalestate_0/un1_timecount_2_sqmuxa_4 ), .Y(
        \scalestate_0/timecount_m1_e_2_2 ));
    IOPAD_IN \ddsclkout_pad/U0/U0  (.PAD(ddsclkout), .Y(
        \ddsclkout_pad/U0/NET1 ));
    AO1 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_45  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[1] )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[2] )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[0] )
        , .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ));
    NOR3A \top_code_0/s_load_RNO_1  (.A(\top_code_0/N_333 ), .B(
        \top_code_0/N_144 ), .C(\top_code_0/N_152 ), .Y(
        \top_code_0/N_302 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[2]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_7_2 ), .Y(
        \timer_top_0/timer_0/timedata_4[2] ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m46_0 ));
    NOR3B \top_code_0/cal_load_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_333 ), .C(\top_code_0/N_155 ), .Y(
        \top_code_0/N_272 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[15]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[15]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_495 ));
    XA1A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_20[10]  (.A(
        \sd_acq_top_0/count[21] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[21]_net_1 ), .C(
        net_27), .Y(\sd_acq_top_0/sd_sacq_coder_0/i_0_0[10] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[20]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[20]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_467 ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_20  (.A(
        \top_code_0_sigtimedata[6] ), .B(
        \ClockManagement_0/long_timer_0/count[6]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_6 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI47Q6[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_6[0] ));
    DFN1E1 \scalestate_0/OPENTIME[5]  (.D(\top_code_0_scaledatain[5] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[5]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[19]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[19]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_507 ));
    OR2A \top_code_0/s_addchoice_1_sqmuxa_0_o2_0  (.A(\xa_c[3] ), .B(
        \top_code_0/N_147 ), .Y(\top_code_0/N_164 ));
    DFN1 \top_code_0/k2  (.D(\top_code_0/k2_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(k2_c));
    NOR2A \DUMP_0/dump_coder_0/para4_4[11]  (.A(
        \top_code_0_dumpdata_0[11] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[11]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[6] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_36  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_42_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_37_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_36_Y ));
    NOR3 \DDS_0/dds_coder_0/i_RNO_0[3]  (.A(\DDS_0/count[3] ), .B(
        \DDS_0/count[1] ), .C(\DDS_0/count[2] ), .Y(
        \DDS_0/dds_coder_0/m8_2 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[0]  (.A(
        \scanstate_0_timecount[0] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_241 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[0]  (.D(
        \PLUSE_0/bri_timer_0/count_e0 ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_8[0] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[9]  (.A(
        \timer_top_0/state_switch_0/N_200 ), .B(
        \timer_top_0/state_switch_0/N_201 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[9] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[9]_net_1 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[14]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_40 ), .Y(
        \timer_top_0/timer_0/timedata_4[14] ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/signal_data_t_0_13  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] ), .Y(
        \Signal_Noise_Acq_0/un1_signal_acq_0[1] ));
    MX2 \nsctrl_choice_0/dumpon_ctr_RNO_0  (.A(scanstate_0_dds_conf), 
        .B(noisestate_0_dumpon_ctr), .S(top_code_0_n_s_ctrl_0), .Y(
        \nsctrl_choice_0/dumpon_ctr_5 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_17[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[13]_net_1 ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_13[0] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[6]  (.D(
        \top_code_0_pd_pluse_data[6] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[6]_net_1 ));
    DFN1 \s_acq_change_0/s_stripnum[4]  (.D(
        \s_acq_change_0/s_stripnum_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[4] ));
    AO1 \state_1ms_0/timecount_RNO_4[13]  (.A(
        \state_1ms_0/S_DUMPTIME[13]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[13] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[13] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[15]_net_1 ));
    DFN1 \plusestate_0/CS[4]  (.D(\plusestate_0/CS_RNO_0[4]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[4]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[3]  (.A(
        \noisestate_0_timecount[3] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_225 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m44 ));
    AOI1 \scalestate_0/CS_RNIVS7S[17]  (.A(\scalestate_0/CS[17]_net_1 )
        , .B(top_code_0_inv_turn), .C(scalestate_0_ne_le), .Y(
        \scalestate_0/N_1265 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[2]_net_1 ));
    DFN1 \s_acq_change_0/s_acqnum[0]  (.D(
        \s_acq_change_0/s_acqnum_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[8] ));
    DFN1E1 \top_code_0/plusedata[15]  (.D(\GPMI_0_dataout[15] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[15] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m179  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_180 ));
    AO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_64  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[2] )
        );
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[6]  (.D(
        \top_code_0_pd_pluse_data[6] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[6]_net_1 ));
    NOR2B \n_acq_change_0/n_rst_n_0  (.A(
        \n_acq_change_0/n_rst_n_5_net_1 ), .B(net_27), .Y(
        \n_acq_change_0/n_rst_n_0_net_1 ));
    DFN1 \s_acq_change_0/s_acqnum[15]  (.D(
        \s_acq_change_0/s_acqnum_RNO[15]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[15] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_60_i ));
    DFN1 \scalestate_0/CS[9]  (.D(\scalestate_0/CS_RNO_0[9]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[9]_net_1 ));
    DFN1E1 \scalestate_0/ACQTIME[14]  (.D(\top_code_0_scaledatain[14] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[14]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_52_i ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[4]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c2 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n4 ));
    DFN1 \scalestate_0/s_acqnum_1[11]  (.D(
        \scalestate_0/s_acqnum_1_RNO[11]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[11] ));
    NOR2B \DUMP_0/off_on_timer_0/count_RNO_0[4]  (.A(
        \DUMP_0/count_2[3] ), .B(\DUMP_0/off_on_timer_0/count_c2 ), .Y(
        \DUMP_0/off_on_timer_0/count_9_0 ));
    NOR3B \DUMP_0/off_on_coder_1/i_RNO_0[1]  (.A(\DUMP_0/count_2[4] ), 
        .B(\DUMP_0/count_2[2] ), .C(\DUMP_0/count_2[3] ), .Y(
        \DUMP_0/off_on_coder_1/i_0_2[1] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m152  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_153 ));
    NOR3B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_RNO[3]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_9_1 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[3] ));
    OR3 \top_code_0/un1_state_1ms_rst_n117_18_i_o2  (.A(\xa_c[6] ), .B(
        \top_code_0/N_137 ), .C(
        \top_code_0/un1_state_1ms_rst_n117_18_i_o2_0_net_1 ), .Y(
        \top_code_0/N_167 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_22  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[3] )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_54  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_60_i ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3_0 ));
    XO1 \PLUSE_0/qq_coder_1/un1_qq_para2_NE_0[0]  (.A(
        \PLUSE_0/count_7[4] ), .B(\PLUSE_0/qq_para2[4] ), .C(
        \PLUSE_0/qq_para2[5] ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_0[0]_net_1 ));
    MX2 \PLUSE_0/bri_coder_0/i[1]/U0  (.A(\PLUSE_0/i_8[1] ), .B(
        \PLUSE_0/bri_coder_0_half ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_coder_0/i[1]/Y ));
    DFN1E1 \plusestate_0/DUMPTIME[0]  (.D(\top_code_0_plusedata[0] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[0]_net_1 ));
    NOR2A \noisestate_0/timecount_1_RNO[14]  (.A(\noisestate_0/N_71 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[14] ));
    MX2 \scanstate_0/timecount_1_RNO_0[2]  (.A(
        \scanstate_0/acqtime[2]_net_1 ), .B(
        \scanstate_0/dectime[2]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_60 ));
    DFN1E1 \top_code_0/scandata[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[3] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIQ7U0A[12]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_17[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_16[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_18[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_i[0] ));
    AO1 \scalestate_0/timecount_ret_60_RNO_2  (.A(
        \scalestate_0/CUTTIME180_TEL[12]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[12] )
        , .Y(\scalestate_0/timecount_20_iv_3[12] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m197  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_198 ));
    MX2B \noisestate_0/timecount_1_RNO[0]  (.A(\noisestate_0/N_57 ), 
        .B(top_code_0_noise_rst_0), .S(\noisestate_0/N_228 ), .Y(
        \noisestate_0/timecount_5[0] ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIV5JJ9[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_14[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_28  (.A(
        \timer_top_0/dataout[7] ), .B(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_28_Y ));
    DFN1 \timer_top_0/state_switch_0/clk_en_scan  (.D(
        \timer_top_0/state_switch_0/clk_en_scan_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(timer_top_0_clk_en_scan));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[11]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[10] )
        , .Y(\DDS_0/dds_state_0/N_325 ));
    MX2 \scanstate_0/timecount_1_RNO_0[4]  (.A(
        \scanstate_0/dectime[4]_net_1 ), .B(
        \scanstate_0/acqtime[4]_net_1 ), .S(\scanstate_0/CS[4]_net_1 ), 
        .Y(\scanstate_0/N_62 ));
    DFN1E1 \scalestate_0/PLUSETIME180[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[13]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[2]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_30  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[5] ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m80  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_79 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_80 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_81 ));
    AO1 \bridge_div_0/dataall_1_I_15  (.A(
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0[0] ), .B(
        \bridge_div_0/DWACT_ADD_CI_0_TMP[0] ), .C(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_1[0] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_1[0] ));
    DFN1 \scalestate_0/s_acqnum_1[0]  (.D(
        \scalestate_0/s_acqnum_1_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[0] ));
    DFN1E1 \scalestate_0/ACQTIME[4]  (.D(\top_code_0_scaledatain[4] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[4]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[9] ));
    DFN1 \DUMP_0/dump_state_0/cs[2]  (.D(
        \DUMP_0/dump_state_0/cs_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[2]_net_1 ));
    DFN1 \scalestate_0/CS[5]  (.D(\scalestate_0/CS_RNO_1[5] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[5]_net_1 ));
    DFN1E1 \top_code_0/noisedata[15]  (.D(\GPMI_0_dataout[15] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[15] ));
    DFN1E1 \top_code_0/scaledatain[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[5] ));
    DFN1E1 \scalestate_0/CUTTIME90[9]  (.D(\top_code_0_scaledatain[9] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[9]_net_1 ));
    DFN1E1 \scalestate_0/timecount[20]  (.D(
        \scalestate_0/timecount_20[20] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(\scalestate_0_timecount[20] ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_2  (.A(
        \scalestate_0/M_NUM[9]_net_1 ), .B(
        \scalestate_0/necount[9]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_2_Y ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[0]  (.D(
        \top_code_0_pd_pluse_data[0] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[0]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[6]_net_1 ));
    NOR2A \scalestate_0/CS_RNO[2]  (.A(top_code_0_scale_rst_3), .B(
        \scalestate_0/CS_srsts_i_0[2] ), .Y(\scalestate_0/CS_RNO_1[2] )
        );
    NOR2B \top_code_0/k2_RNO_3  (.A(\xa_c[1] ), .B(\xa_c[5] ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_2 ));
    OA1B \syn_md_module_1/syn_md_0/count_RNO[3]  (.A(
        \syn_md_module_1/syn_md_0/N_23_1 ), .B(
        \syn_md_module_1/syn_md_0/N_22 ), .C(
        \syn_md_module_1/syn_md_0/N_50 ), .Y(
        \syn_md_module_1/syn_md_0/count_RNO[3]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[7]_net_1 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIS7HQ[15]  (
        .A(\pd_pluse_top_0/count[15] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[15]_net_1 ), 
        .C(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_14[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_0[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m141  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_138 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_141 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_142 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNITB6T[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[10]_net_1 ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_10[0] ));
    NOR3C \scalestate_0/timecount_ret_50_RNO_1  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[17]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[17] ));
    NOR3C \scalestate_0/M_NUM_1_sqmuxa_0_a2  (.A(
        \top_code_0_scalechoice_0[0] ), .B(\scalestate_0/N_61 ), .C(
        \scalestate_0/N_64 ), .Y(\scalestate_0/M_NUM_1_sqmuxa ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_40_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m42_5 ));
    OR2B \scalestate_0/bb_ch_RNO_1  (.A(\scalestate_0/un1_CS_20 ), .B(
        timer_top_0_clk_en_scale), .Y(\scalestate_0/N_1177 ));
    NOR2A \state_1ms_0/M_DUMPTIME_1_sqmuxa_0_a2_0  (.A(
        \state_1ms_0/N_16 ), .B(\top_code_0_state_1ms_lc[2] ), .Y(
        \state_1ms_0/N_17 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[26]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[26]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_471 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[5]  (.D(
        \top_code_0_bri_datain[15] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/qq_para3[5] ));
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en  (.A(
        n_acq_change_0_n_acq_start), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0_en ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en_net_1 ));
    NOR2B \PLUSE_0/bri_timer_0/count_RNILIEB[5]  (.A(
        \PLUSE_0/bri_timer_0/count_c4 ), .B(\PLUSE_0/count_2[5] ), .Y(
        \PLUSE_0/bri_timer_0/count_c5 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_38  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_38_Y ));
    OR3 \DUMP_0/dump_coder_0/para2_RNIGTH12[2]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_3[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_3_4[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_3_NE_3[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_7[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[8]_net_1 ));
    AOI1A \PLUSE_0/bri_coder_0/half_0_I_13  (.A(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[3] ), .B(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[4] ), .C(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[5] ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[0] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_10  (.A(
        \timer_top_0/dataout[4] ), .B(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_10_Y ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[14]  (.D(
        \top_code_0_state_1ms_data[14] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[14]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[11]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNICLLJ[1]  (.A(
        \DUMP_0/dump_coder_0/para5[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_0[0] ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[17]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[17]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[6]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[6]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[6] ));
    AO1 \DUMP_0/dump_state_0/off_start_RNO  (.A(
        \DUMP_0/dump_state_0/N_176 ), .B(\DUMP_0/dump_state_0/cs4 ), 
        .C(\DUMP_0/dump_state_0/cs_nsss[6] ), .Y(
        \DUMP_0/dump_state_0/off_start_RNO_net_1 ));
    AND3 \scalestate_0/necount_inc_0/FND2_9_inst  (.A(
        \scalestate_0/necount_inc_0/inc_12_net ), .B(
        \scalestate_0/necount_inc_0/inc_5_net ), .C(
        \scalestate_0/necount_inc_0/inc_10_net ), .Y(
        \scalestate_0/necount_inc_0/Rcout_10_net ));
    NOR2B \scalestate_0/bb_ch_RNO  (.A(\scalestate_0/N_729 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/bb_ch_RNO_net_1 ));
    NOR3A \top_code_0/scan_start_ret_2_RNO  (.A(
        \top_code_0/un1_xa_10_2 ), .B(\top_code_0/N_144 ), .C(
        \top_code_0/N_165 ), .Y(\top_code_0/un1_xa_10 ));
    MX2 \top_code_0/relay_close_RNO_0[3]  (.A(\relay_close_c[3] ), .B(
        \GPMI_0_dataout[3] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_822 ));
    OA1C \top_code_0/pluse_scale_RNO_0  (.A(\xa_c[1] ), .B(
        \top_code_0/N_176 ), .C(top_code_0_pluse_scale), .Y(
        \top_code_0/N_295 ));
    DFN1E1 \scalestate_0/ACQTIME[10]  (.D(\top_code_0_scaledatain[10] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[10]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_66_i ));
    IOPAD_IN \xa_pad[10]/U0/U0  (.PAD(xa[10]), .Y(\xa_pad[10]/U0/NET1 )
        );
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_56_i ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[3]  (.A(
        \DUMP_0/dump_timer_0/count_c2 ), .B(\DUMP_0/count_1[3] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n3 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[1]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[1]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_280 ));
    NOR2B \sd_acq_top_0/sd_sacq_state_0/cs_RNILI5E[9]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[9]_net_1 ), .B(
        \sd_acq_top_0/i_0[7] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_232 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_83  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_83_Y ));
    IOPAD_IN \ADC_pad[2]/U0/U0  (.PAD(ADC[2]), .Y(\ADC_pad[2]/U0/NET1 )
        );
    DFN1 \DUMP_0/off_on_state_0/state_over  (.D(
        \DUMP_0/off_on_state_0/N_9 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/off_on_state_0_state_over ));
    MX2 \noisestate_0/timecount_1_RNO[2]  (.A(\noisestate_0/N_59 ), .B(
        \noisestate_0/timecount_cnst[2] ), .S(\noisestate_0/N_228 ), 
        .Y(\noisestate_0/timecount_5[2] ));
    NOR2B \scalestate_0/strippluse_RNO[0]  (.A(\scalestate_0/N_559 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[0]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[8]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[8] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[8]_net_1 )
        );
    DFN1E1 \top_code_0/s_periodnum[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_periodnum_1_sqmuxa ), .Q(
        \top_code_0_s_periodnum[3] ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_11  (.A(
        \timer_top_0/dataout[10] ), .B(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_12_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_11_Y ));
    OR2A \top_code_0/un1_xa_30_0_o2_0  (.A(\top_code_0/N_13 ), .B(
        \top_code_0/N_127 ), .Y(\top_code_0/un1_xa_30_0_o2_0_net_1 ));
    DFN1E1 \top_code_0/dumpdata[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[9] ));
    MX2 \scalestate_0/long_opentime_RNO_0  (.A(
        \scalestate_0/necount_LE_M_net_1 ), .B(
        scalestate_0_long_opentime), .S(\scalestate_0/N_1163 ), .Y(
        \scalestate_0/N_743 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIADQ6[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_9[0] ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[5]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_2[5] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[5]_net_1 )
        );
    MX2 \scanstate_0/timecount_1_RNO[4]  (.A(\scanstate_0/N_62 ), .B(
        \scanstate_0/timecount_cnst[4] ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[4] ));
    NOR3C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[4]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/i_1[3] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs[3]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[4] ));
    XOR2 \bridge_div_0/count_5_I_5  (.A(
        \bridge_div_0/count_RNIEMOM7[0]_net_1 ), .B(
        \bridge_div_0/count_RNIFNOM7[1]_net_1 ), .Y(
        \bridge_div_0/count_5[1] ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[3]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[3] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[3] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[8]  (.A(\scalestate_0/N_456 ), 
        .B(\scalestate_0/ACQECHO_NUM[8]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[8] ));
    AND2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_21  
        (.A(\s_acq_change_0_s_stripnum[6] ), .B(
        \s_acq_change_0_s_stripnum[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[3] )
        );
    NOR2B \DUMP_0/dump_coder_0/i_RNO[2]  (.A(
        state1ms_choice_0_bri_cycle), .B(state1ms_choice_0_reset_out), 
        .Y(\DUMP_0/dump_coder_0/i_RNO_0[2] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[7]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[7] ));
    OR2B \scalestate_0/CS_RNIKLDI[6]  (.A(\scalestate_0/CS[6]_net_1 ), 
        .B(top_code_0_scale_rst), .Y(\scalestate_0/N_1069 ));
    NOR2A \top_code_0/change_1_sqmuxa_0_a2_0  (.A(net_27), .B(
        \top_code_0/N_148 ), .Y(\top_code_0/N_331 ));
    AO1 \timer_top_0/state_switch_0/dataout_RNO[19]  (.A(
        \state_1ms_0_timecount[19] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .C(
        \timer_top_0/state_switch_0/N_272 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[19]_net_1 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[9]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[9] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[9]_net_1 ));
    AO1A \scalestate_0/timecount_ret_70_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/S_DUMPTIME[15]_net_1 ), .C(
        \scalestate_0/timecount_20_iv_1[15] ), .Y(
        \scalestate_0/timecount_20_iv_6[15] ));
    NOR3B \DDS_0/dds_state_0/data_RNO  (.A(
        \DDS_0/dds_state_0/para[0]_net_1 ), .B(
        \DDS_0/dds_state_0/N_223 ), .C(\DDS_0/dds_state_0/N_531 ), .Y(
        \DDS_0/dds_state_0/N_21 ));
    DFN1 \s_acq_change_0/s_acqnum[2]  (.D(
        \s_acq_change_0/s_acqnum_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[2] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[8]  (.D(
        \top_code_0_state_1ms_data[8] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[8]_net_1 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3_I_7  (
        .A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIKJJB2[2]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[2] ));
    DFN1E1 \scalestate_0/timecount_ret_87  (.D(
        \scalestate_0/timecount_20_iv_2[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_2_reto[10] ));
    NOR3C \DUMP_0/dump_coder_0/i_RNO[3]  (.A(
        \DUMP_0/dump_coder_0/N_19 ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] ), .C(
        \DUMP_0/dump_coder_0/i_0_0_a2_12[3] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO_0[3]_net_1 ));
    IOIN_IB \ADC_pad[9]/U0/U1  (.YIN(\ADC_pad[9]/U0/NET1 ), .Y(
        \ADC_c[9] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m88  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_87 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_88 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_89 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[13]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[12] )
        , .Y(\DDS_0/dds_state_0/N_334 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[4]  (.A(
        \plusestate_0_timecount[4] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_224 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m194  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_195 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n2 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2]/Y ));
    NOR2 \scalestate_0/CS_RNIPB6E[18]  (.A(\scalestate_0/CS[18]_net_1 )
        , .B(\scalestate_0/N_1201 ), .Y(
        \scalestate_0/un1_CS6_39_i_a2_0 ));
    DFN1E0 \DDS_0/dds_state_0/para[13]  (.D(\DDS_0/dds_state_0/N_118 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[13]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[0]  (.A(
        \plusestate_0_timecount[0] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_244 ));
    IOPAD_TRI \relay_close_pad[9]/U0/U0  (.D(
        \relay_close_pad[9]/U0/NET1 ), .E(\relay_close_pad[9]/U0/NET2 )
        , .PAD(relay_close[9]));
    NOR2A \GPMI_0/tri_state_0/dataout_1_11  (.A(\xd_in[3] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[3] ));
    NOR3A \ClockManagement_0/long_timer_0/timeup_RNO_12  (.A(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_4 ), .B(
        \ClockManagement_0/long_timer_0/clear_n4_1 ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_2 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_10 ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa_0_a2_0  
        (.A(top_code_0_sd_sacq_load), .B(
        \top_code_0_sd_sacq_choice[2] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_0  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I10_un1_CO1 ), 
        .B(\s_acq_change_0_s_stripnum[11] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_11 )
        );
    AO1A \scalestate_0/timecount_ret_40_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[2]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[2] ), .Y(
        \scalestate_0/timecount_20_iv_1[2] ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[17]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_49 ), .Y(
        \timer_top_0/timer_0/timedata_4[17] ));
    DFN1 \DDS_0/dds_coder_0/i[3]  (.D(
        \DDS_0/dds_coder_0/i_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/i[3] ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_32  (.A(
        \timer_top_0/timer_0/N_12 ), .B(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .Y(
        \timer_top_0/timer_0/I_32_2 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[15]_net_1 ));
    NOR2B \PLUSE_0/qq_timer_1/count_RNO_0[4]  (.A(\PLUSE_0/count_7[3] )
        , .B(\PLUSE_0/qq_timer_1/count_c2 ), .Y(
        \PLUSE_0/qq_timer_1/count_9_0 ));
    OR3 \scalestate_0/timecount_ret_71_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[15] ), .B(
        \scalestate_0/OPENTIME_TEL_m[15] ), .C(
        \scalestate_0/timecount_20_iv_4[15] ), .Y(
        \scalestate_0/timecount_20_iv_8[15] ));
    DFN1E1 \noisestate_0/dectime[1]  (.D(\top_code_0_noisedata[1] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[1]_net_1 ));
    DFN1E1 \top_code_0/pluse_scale  (.D(\top_code_0/N_88 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pluse_scale));
    DFN1E1 \top_code_0/pd_pluse_data[9]  (.D(\GPMI_0_dataout[9] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[9] ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[3]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[3] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/en1 ));
    NOR3A \sd_acq_top_0/sd_sacq_coder_0/i_RNO[7]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[7] ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[4]  (.A(
        \top_code_0_dumpdata_0[4] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[4]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[4]  (.A(
        \noisestate_0_timecount[4] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_220 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m39  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_40 ));
    AO1C \plusestate_0/CS_RNO_0[6]  (.A(\plusestate_0/CS[5]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst), .Y(
        \plusestate_0/CS_srsts_i_0[6] ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNICME74[7]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_3[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_2[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_8[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_12[0] ));
    AO1B \scalestate_0/reset_out_RNO_2  (.A(
        \scalestate_0/un1_CS6_39_i_a3_1 ), .B(\scalestate_0/N_1304 ), 
        .C(timer_top_0_clk_en_scale), .Y(\scalestate_0/N_1189 ));
    OAI1 \noisestate_0/CS_RNIOJ68[2]  (.A(\noisestate_0/CS[4]_net_1 ), 
        .B(\noisestate_0/CS[2]_net_1 ), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/N_228 ));
    DFN1 \DUMP_0/off_on_state_1/state_over  (.D(
        \DUMP_0/off_on_state_1/N_9 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/off_on_state_1_state_over ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i10_mux ));
    DFN1 \scalestate_0/bb_ch  (.D(\scalestate_0/bb_ch_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(net_51));
    NOR2B \PLUSE_0/qq_timer_1/count_RNIF2RU[1]  (.A(
        \PLUSE_0/count_7[1] ), .B(\PLUSE_0/count_7[0] ), .Y(
        \PLUSE_0/qq_timer_1/count_c1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m149  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_148 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_149 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_150 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i14_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_106  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_106_Y ));
    DFN1E1 \scalestate_0/timecount_ret_47  (.D(
        \scalestate_0/timecount_20_0_iv_4[16] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_4_reto[16] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[9]  (.A(
        \scalestate_0/ACQ180_NUM[9]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[9]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_457 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[1]  (.D(
        \ClockManagement_0/long_timer_0/count_n1 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[1]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[16]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[16]_net_1 ));
    DFN1E1 \scalestate_0/DUMPTIME[5]  (.D(\top_code_0_scaledatain[5] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[5]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[0]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[0] ));
    NOR2B \scalestate_0/timecount_ret_28_RNO_5  (.A(
        \scalestate_0/CUTTIME180[1]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[1] ));
    NOR3C \CAL_0/cal_div_0/count_RNO[1]  (.A(net_33_0), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(\CAL_0/cal_div_0/I_5 ), 
        .Y(\CAL_0/cal_div_0/count_5[1] ));
    NOR2B \top_code_0/relay_close_RNO[8]  (.A(\top_code_0/N_827 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[8]_net_1 ));
    RAM512X18 #( .MEMORYFILE("RAM_R5C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R5C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_5_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_5_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_0_net ));
    NOR2B \DUMP_0/dump_coder_0/i_RNO[0]  (.A(
        state1ms_choice_0_dump_start), .B(state1ms_choice_0_reset_out), 
        .Y(\DUMP_0/dump_coder_0/i_RNO_0[0] ));
    DFN1 \DUMP_ON_0/off_on_state_0/cs[1]  (.D(
        \DUMP_ON_0/off_on_state_0/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/off_on_state_0/cs[1]_net_1 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_9  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_3_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_4_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_10_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_9_Y ));
    NOR3A \top_code_0/k2_RNO_4  (.A(\xa_c[7] ), .B(\xa_c[18] ), .C(
        \top_code_0/N_127 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_1 ));
    NOR3C \PLUSE_0/qq_timer_1/count_0_sqmuxa  (.A(
        \PLUSE_0/qq_state_1_stateover ), .B(\PLUSE_0/down ), .C(
        bri_dump_sw_0_reset_out), .Y(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[3]  (.A(
        \top_code_0_dumpdata_0[3] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[3]_net_1 ));
    OR2A \scalestate_0/necount_cmp_0/OR2A_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/M_NUM[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_3_Y ));
    DFN1E1 \top_code_0/scaleddsdiv[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[4] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]  (.D(
        \top_code_0_n_acqnum_2[5] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[6]  (.D(
        \top_code_0_pd_pluse_data[6] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[6]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n1 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1]/Y ));
    DFN1 \top_code_0/state_1ms_start_ret  (.D(
        top_code_0_state_1ms_start), .CLK(GLA_net_1), .Q(
        \top_code_0/top_code_0_state_1ms_start_reto ));
    DFN1E1 \top_code_0/scandata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[5] ));
    DFN1E1 \scalestate_0/timecount_ret_82  (.D(
        \scalestate_0/timecount_20_iv_6[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[4] ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIGLFH[4]  (.A(
        \DUMP_0/dump_coder_0/para3[4]_net_1 ), .B(\DUMP_0/count_1[4] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_4[0] ));
    DFN1E1 \top_code_0/bridge_load_0  (.D(\top_code_0/N_62 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_bridge_load_0));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[6]  (.A(
        \noisestate_0_timecount[6] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_210 ));
    DFN1E1 \noisestate_0/acqtime[1]  (.D(\top_code_0_noisedata[1] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[1]_net_1 ));
    NOR2B \top_code_0/state_1ms_start_ret_1_RNINE421  (.A(
        \top_code_0/N_796_reto ), .B(\top_code_0/net_27_reto ), .Y(
        top_code_0_scan_start));
    NOR2B \topctrlchange_0/rt_sw_RNO  (.A(\topctrlchange_0/N_12 ), .B(
        net_27), .Y(\topctrlchange_0/rt_sw_RNO_4 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_3_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[8]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m55  
        (.A(\s_acq_change_0_s_stripnum[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[4]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i6_mux ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_56_i ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIJQ983[8]  (.A(
        \DUMP_0/dump_timer_0/count_c7 ), .B(\DUMP_0/count[8] ), .Y(
        \DUMP_0/dump_timer_0/count_c8 ));
    DFN1E1 \scalestate_0/OPENTIME[4]  (.D(\top_code_0_scaledatain[4] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[4]_net_1 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/FND2_9_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_12_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net )
        , .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_10_net ));
    DFN1 \state_1ms_0/soft_dump  (.D(\state_1ms_0/soft_dump_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(state_1ms_0_soft_dump));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[6]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n6 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[6] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[18]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[18]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[4]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_90  (.D(
        \scalestate_0/timecount_20_iv_2[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_2_reto[8] ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[3]_net_1 ));
    MX2 \scalestate_0/necount_RNO_0[3]  (.A(\scalestate_0/necount1[3] )
        , .B(\scalestate_0/necount[3]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_733 ));
    NOR2B \dds_change_0/dds_conf_RNO_2  (.A(scalestate_0_dds_conf), .B(
        \top_code_0_change[0] ), .Y(\dds_change_0/dds_confin2_m ));
    DFN1P0 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/entop  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/entop_RNO_net_1 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .PRE(
        s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop ));
    DFN1E1 \scalestate_0/timecount_ret_14  (.D(
        \scalestate_0/timecount_20_iv_7[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[9] ));
    MX2B \PLUSE_0/bri_state_0/cs_RNO[8]  (.A(
        \PLUSE_0/bri_state_0/cs[8]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[7] ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_1[8] ));
    NOR3A \DDS_0/dds_state_0/data_RNO_0  (.A(\DDS_0/dds_state_0/N_224 )
        , .B(\DDS_0/dds_state_0/cs[4]_net_1 ), .C(
        \DDS_0/dds_state_0/cs[5]_net_1 ), .Y(\DDS_0/dds_state_0/N_531 )
        );
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[17]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[17]_net_1 ));
    XOR2 \bridge_div_0/datahalf_RNI85JN[1]  (.A(
        \bridge_div_0/datahalf[1]_net_1 ), .B(
        \bridge_div_0/count[1]_net_1 ), .Y(
        \bridge_div_0/clear1_n17_1[0] ));
    NOR2B \scalestate_0/timecount_ret_60_RNO_0  (.A(
        \scalestate_0/CUTTIME180[12]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[12] ));
    MX2 \noisestate_0/timecount_1_RNO_0[2]  (.A(
        \noisestate_0/acqtime[2]_net_1 ), .B(
        \noisestate_0/dectime[2]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_59 ));
    NOR3C \DUMP_0/off_on_coder_1/i_RNO[1]  (.A(
        \DUMP_0/off_on_coder_1/i_0_2[1] ), .B(
        \DUMP_0/off_on_coder_1/i_0_1[1] ), .C(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_coder_1/i_RNO_1[1]_net_1 ));
    DFN1E1 \scanstate_0/dectime[13]  (.D(\top_code_0_scandata[13] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[13]_net_1 ));
    NOR2A \PLUSE_0/qq_coder_0/i_RNO[3]  (.A(bri_dump_sw_0_reset_out), 
        .B(\PLUSE_0/qq_coder_0/i_reg10_NE[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/i_RNO_2[3] ));
    NOR2B \top_code_0/relay_on_RNO[1]  (.A(\top_code_0/N_810 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[1]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[14]  (.D(\GPMI_0_dataout[14] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[14] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIBGT7[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_9[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[4] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m43 ));
    OR2B \noisestate_0/CS_RNIRL68[1]  (.A(\noisestate_0/CS[1]_net_1 ), 
        .B(top_code_0_noise_rst), .Y(\noisestate_0/N_193 ));
    NOR3A \DUMP_0/dump_state_0/cs_RNO[5]  (.A(
        \DUMP_0/dump_state_0/cs4 ), .B(\DUMP_0/dump_state_0/N_193 ), 
        .C(\DUMP_0/dump_state_0/cs_RNO_1[5]_net_1 ), .Y(
        \DUMP_0/dump_state_0/cs_RNO_0[5]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m42_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[17] ));
    DFN1 \timer_top_0/timer_0/timedata[10]  (.D(
        \timer_top_0/timer_0/timedata_4[10] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[10]_net_1 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_10_RNO_1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N160 ), 
        .B(\s_acq_change_0_s_stripnum[8] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_8 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[1] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI6D09[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[11]_net_1 ));
    NOR2B \topctrlchange_0/soft_dump_6_iv_RNO  (.A(scalestate_0_soft_d)
        , .B(\top_code_0_change[0] ), .Y(\topctrlchange_0/s_dumpin2_m )
        );
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[14]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[14] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_0[14] ));
    DFN1 \scalestate_0/dump_start  (.D(
        \scalestate_0/dump_start_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_dump_start));
    XOR2 \PLUSE_0/bri_timer_0/count_RNO[1]  (.A(\PLUSE_0/count_8[0] ), 
        .B(\PLUSE_0/count_8[1] ), .Y(\PLUSE_0/bri_timer_0/count_n1 ));
    AND3B \top_code_0/sd_sacq_data_1_sqmuxa_0_a2  (.A(
        \top_code_0/N_147 ), .B(\top_code_0/N_163 ), .C(
        \top_code_0/N_331 ), .Y(\top_code_0/sd_sacq_data_1_sqmuxa ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[6]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIFGET[11]  (.A(
        \DUMP_0/dump_coder_0/para6[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_11[0] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[1]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m47_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[4] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_41_i ));
    NOR2B \scalestate_0/CS_RNO[17]  (.A(\scalestate_0/N_1230 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[17]_net_1 ));
    DFN1 \top_code_0/pluse_str  (.D(\top_code_0/pluse_str_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(top_code_0_pluse_str));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_9  (.A(
        \timer_top_0/dataout[14] ), .B(
        \timer_top_0/timer_0/timedata[14]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_9_Y ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[9]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[9] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[9] ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIHOII[4]  (.A(
        \DUMP_0/dump_coder_0/para4[4]_net_1 ), .B(\DUMP_0/count_1[4] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_4[0] ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_38  (.A(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[8] ));
    AND2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/FND2_8_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_12_net ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m90  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_91 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1  (.A(\xd_in[15] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[15] ));
    NOR2B \DUMP_0/off_on_coder_1/i_RNO[0]  (.A(
        \DUMP_0/dump_state_0_off_start ), .B(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_coder_1/i_RNO_1[0] ));
    IOPAD_IN \tri_ctrl_pad/U0/U0  (.PAD(tri_ctrl), .Y(
        \tri_ctrl_pad/U0/NET1 ));
    XO1 \DUMP_0/dump_coder_0/para6_RNIC3I91[6]  (.A(
        \DUMP_0/count_0[6] ), .B(\DUMP_0/dump_coder_0/para6[6]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/i_reg16_5[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_1[0] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_50  (.A(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[12] ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[13]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[13] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[13] ));
    OR2 \scalestate_0/CS_RNII6HJ[2]  (.A(\scalestate_0/CS[2]_net_1 ), 
        .B(\scalestate_0/CS[8]_net_1 ), .Y(\scalestate_0/N_1203 ));
    NOR2A \top_code_0/un1_state_1ms_rst_n117_i_a2_0  (.A(\xa_c[1] ), 
        .B(\top_code_0/N_150 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_i_a2_0_net_1 ));
    MX2 \PLUSE_0/bri_coder_0/i[2]/U0  (.A(\PLUSE_0/i_3[2] ), .B(
        bri_dump_sw_0_phase_ctr), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_coder_0/i[2]/Y ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[1]  (.A(
        \timer_top_0/state_switch_0/N_235 ), .B(
        \timer_top_0/state_switch_0/N_236 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[1] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[1]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_67  (.D(
        \scalestate_0/timecount_20_iv_6[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[14] ));
    MX2 \scalestate_0/strippluse_RNO_0[1]  (.A(
        \scalestate_0/strippluse_6[1] ), .B(
        \scalestate_0_strippluse[1] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_560 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[10]  (.D(
        \DUMP_0/dump_coder_0/para2_4[10]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[10]_net_1 ));
    NOR2 \DDS_0/dds_state_0/para_9_i_0_a2_5[22]  (.A(\DDS_0/i[0] ), .B(
        top_code_0_dds_load), .Y(\DDS_0/dds_state_0/N_535 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[14]_net_1 ));
    DFN1 \DUMP_0/dump_coder_0/i[8]  (.D(
        \DUMP_0/dump_coder_0/i_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i[8] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[20]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[20]_net_1 ));
    DFN1 \scanstate_0/CS[5]  (.D(\scanstate_0/CS_RNO_2[5] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[5]_net_1 ));
    XOR2 \bridge_div_0/dataall_RNI6UNO[1]  (.A(
        \bridge_div_0/dataall[1]_net_1 ), .B(
        \bridge_div_0/count[1]_net_1 ), .Y(
        \bridge_div_0/un1_count_1_0[0] ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[4]_net_1 ));
    AO1C \PLUSE_0/bri_coder_0/half_0_I_20  (.A(\PLUSE_0/half_para[2] ), 
        .B(\PLUSE_0/count_8[2] ), .C(\PLUSE_0/bri_coder_0/N_2 ), .Y(
        \PLUSE_0/bri_coder_0/N_8 ));
    DFN1 \ClockManagement_0/clk_10k_0/count[1]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[1] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[1]_net_1 ));
    NOR3 \top_code_0/dds_choice_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_164 ), .Y(
        \top_code_0/N_274 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[10]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n10 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[6]  (.A(
        \sd_acq_top_0/i_2[4] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_219 ));
    AND3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_8  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3 ));
    MX2 \top_code_0/relay_on_RNO_0[0]  (.A(\relay_on_c[0] ), .B(
        \GPMI_0_dataout[0] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_809 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_1_inst  (.A(
        \sd_acq_top_0/count_10[0] ), .B(\sd_acq_top_0/count_10[1] ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/count1[1] ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[7]  (.D(
        \DUMP_0/dump_coder_0/para4_4[7]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[7]_net_1 ));
    RAM512X18 #( .MEMORYFILE("RAM_R8C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R8C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_8_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_8_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_0_net ));
    DFN1E1 \scanstate_0/timecount_1[11]  (.D(
        \scanstate_0/timecount_5[11] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[11] ));
    NOR3B \PLUSE_0/qq_coder_0/i_RNO[2]  (.A(bri_dump_sw_0_reset_out), 
        .B(\PLUSE_0/qq_coder_0/i_reg10_NE[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_0/un1_qq_para2_i[0] ), .Y(
        \PLUSE_0/qq_coder_0/i_RNO_2[2] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m47_1 ));
    OR2A \scalestate_0/CS6_0_o2  (.A(top_code_0_scale_rst_5), .B(
        timer_top_0_clk_en_scale), .Y(\scalestate_0/N_1196 ));
    XA1C \DUMP_0/dump_coder_0/i_RNO_8[3]  (.A(\DUMP_0/count_1[0] ), .B(
        \DUMP_0/dump_coder_0/para1[0]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_1[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_1[3] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[5]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[5] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_0_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_165_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_34_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_0_inst ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_2_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/count_10[3] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[3] ));
    AO1 \scalestate_0/timecount_ret_50_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[17]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[17] ), .Y(
        \scalestate_0/timecount_20_0_iv_2[17] ));
    DFN1E1 \scalestate_0/timecount_ret_50  (.D(
        \scalestate_0/timecount_20_0_iv_4[17] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_4_reto[17] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[1] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[26]  (.D(
        \top_code_0_dds_configdata[9] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[26]_net_1 ));
    DFN1 \timer_top_0/timer_0/timedata[11]  (.D(
        \timer_top_0/timer_0/timedata_4[11] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[11]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_7_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_116_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_143_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_7_inst ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNIVADS[2]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c2 ));
    DFN1E1 \noisestate_0/dectime[11]  (.D(\top_code_0_noisedata[11] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[11]_net_1 ));
    DFN1 \scalestate_0/CS[7]  (.D(\scalestate_0/CS_RNO_1[7] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[7]_net_1 ));
    IOPAD_TRI \syn_md_tmp_pad/U0/U0  (.D(\syn_md_tmp_pad/U0/NET1 ), .E(
        \syn_md_tmp_pad/U0/NET2 ), .PAD(syn_md_tmp));
    DFN1E1 \scalestate_0/CUTTIMEI90[21]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[21]_net_1 )
        );
    DFN1C0 \PLUSE_0/bri_state_0/cs[3]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[3] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[3]_net_1 ));
    IOTRI_OB_EB \relay_close_pad[2]/U0/U1  (.D(\relay_close_c[2] ), .E(
        VCC), .DOUT(\relay_close_pad[2]/U0/NET1 ), .EOUT(
        \relay_close_pad[2]/U0/NET2 ));
    NOR2 \scanstate_0/sw_acq2_RNO_1  (.A(\scanstate_0/CS[3]_net_1 ), 
        .B(\scanstate_0/CS[4]_net_1 ), .Y(\scanstate_0/N_238 ));
    NOR2B \state_1ms_0/timecount_RNO_3[11]  (.A(
        \state_1ms_0/CUTTIME[11]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[11] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n7 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        );
    MX2 \nsctrl_choice_0/rt_sw_RNO_0  (.A(scanstate_0_rt_sw), .B(
        noisestate_0_rt_sw), .S(top_code_0_n_s_ctrl_0), .Y(
        \nsctrl_choice_0/rt_sw_5 ));
    OA1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIKJJB2[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIKJJB2[2]_net_1 )
        );
    OR2 \top_code_0/un1_state_1ms_rst_n117_3_4_i_0_o3  (.A(\xa_c[9] ), 
        .B(\xa_c[8] ), .Y(\top_code_0/N_127 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNICCFQ1[21]  (.A(
        \sd_acq_top_0/count[21] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[21]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_17[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_0[0] ));
    DFN1E1 \top_code_0/scalechoice[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0[3] ));
    OA1B \scanstate_0/CS_RNO[7]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[7]_net_1 ), .C(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Y(
        \scanstate_0/CS_RNO_2[7] ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[13]  
        (.D(\s_acq_change_0_s_acqnum[13] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[13]_net_1 )
        );
    DFN1E1 \top_code_0/sd_sacq_data[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[11] ));
    IOPAD_TRI \soft_dump_pad/U0/U0  (.D(\soft_dump_pad/U0/NET1 ), .E(
        \soft_dump_pad/U0/NET2 ), .PAD(soft_dump));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[13]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[13] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count[13] ));
    AO1D \timer_top_0/timer_0/Timer_Cmp_0/AO1D_0  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_4_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_5_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_8_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1D_0_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_74  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_74_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[30]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[30]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_514 ));
    DFN1E1 \top_code_0/s_acqnum[12]  (.D(\GPMI_0_dataout[12] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[12] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_6  (.A(
        \timer_top_0/dataout[10] ), .B(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_6_Y ));
    NOR3 \top_code_0/nstatechoice_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_164 ), .Y(
        \top_code_0/N_286 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m227  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_228 ));
    DFN1E1 \state_1ms_0/CUTTIME[4]  (.D(\top_code_0_state_1ms_data[4] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[4]_net_1 ));
    NOR2B \ClockManagement_0/clk_div500_0/un1_count_1_I_42  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] ), 
        .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_1_1[0] )
        , .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_11[0] ));
    OR2A \plusestate_0/CS_RNI268Q[6]  (.A(top_code_0_pluse_rst), .B(
        \plusestate_0/N_302 ), .Y(\plusestate_0/un1_sw_acq1_2_sqmuxa ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[5]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[5]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_321 ));
    MX2 \plusestate_0/timecount_1_RNO_0[1]  (.A(
        \plusestate_0/DUMPTIME[1]_net_1 ), .B(
        \plusestate_0/PLUSETIME[1]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_72 ));
    NOR2B \DUMP_0/dump_state_0/cs_RNO[7]  (.A(
        \DUMP_0/dump_state_0/N_168 ), .B(\DUMP_0/dump_state_0/cs4 ), 
        .Y(\DUMP_0/dump_state_0/cs_nsss[7] ));
    DFN1E1 \scalestate_0/timecount_ret_62  (.D(
        \scalestate_0/timecount_20_iv_8[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[12] ));
    OR3 \PLUSE_0/qq_coder_0/un1_qq_para2_NE[0]  (.A(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_1[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_0[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_i[0] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[14]  (.A(
        \timer_top_0/state_switch_0/N_262 ), .B(
        \timer_top_0/state_switch_0/N_264 ), .C(
        \timer_top_0/state_switch_0/N_263 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[14] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[0]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_i ));
    NOR3A \top_code_0/k1_RNO_2  (.A(
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_2 ), .B(
        \top_code_0/N_127 ), .C(\xa_c[4] ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_4 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_18  (.A(
        \timer_top_0/dataout[5] ), .B(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_18_Y ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m62  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[0] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_63 ));
    NOR2B \PLUSE_0/bri_state_0/cs_RNO_6[3]  (.A(
        \PLUSE_0/bri_state_0/cs_i_0[12] ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[6] ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_1 ));
    NOR3C \scalestate_0/PLUSETIME180_1_sqmuxa_0_a2  (.A(
        \top_code_0_scalechoice_0[0] ), .B(\scalestate_0/N_61 ), .C(
        \scalestate_0/N_62 ), .Y(\scalestate_0/PLUSETIME180_1_sqmuxa ));
    DFN1 \s_acq_change_0/s_stripnum[11]  (.D(
        \s_acq_change_0/s_stripnum_RNO[11]_net_1 ), .CLK(GLA_net_1), 
        .Q(\s_acq_change_0_s_stripnum[11] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m98  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_99 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[14]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[14]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_463 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[1]  (.D(
        \top_code_0_bri_datain[11] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para3[1] ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNINQCG[8]  (.A(
        \DUMP_0/dump_coder_0/para2[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_8[0] ));
    NOR2B \noisestate_0/dumpoff_ctr_RNO  (.A(\noisestate_0/N_112 ), .B(
        top_code_0_noise_rst), .Y(
        \noisestate_0/dumpoff_ctr_RNO_0_net_1 ));
    OR2 \scalestate_0/reset_out_RNO_3  (.A(\scalestate_0/CS[6]_net_1 ), 
        .B(\scalestate_0/N_1212 ), .Y(\scalestate_0/un1_CS_44_i_0 ));
    NOR2A \plusestate_0/pluse_acq_RNO_1  (.A(\plusestate_0/N_301 ), .B(
        \plusestate_0/CS[9]_net_1 ), .Y(\plusestate_0/N_305 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[9]_net_1 ));
    AND3 \scalestate_0/necount_inc_0/AND2b_9_inst  (.A(
        \scalestate_0/necount[0]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .C(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/incb_2_net ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[18]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[18] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[18] ));
    NOR2 \state_1ms_0/pluse_start_RNO_1  (.A(\state_1ms_0/CS[4]_net_1 )
        , .B(\state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/N_254 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[7]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[7] ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[5]  (.D(
        \top_code_0_cal_data[5] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[5] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_9_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_50_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_32_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_9_inst ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_47  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_47_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_101  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_101_Y ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[21]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[21] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[21] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[25]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[25]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_307 ));
    OA1C \top_code_0/n_load_RNO  (.A(\top_code_0/N_201 ), .B(
        top_code_0_n_load), .C(\top_code_0/N_280 ), .Y(
        \top_code_0/N_72 ));
    MX2 \state1ms_choice_0/rt_sw_RNO  (.A(rt_sw_net_0), .B(
        state_1ms_0_rt_sw), .S(top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/rt_sw_4 ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_24  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[4]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[0] )
        );
    DFN1E1 \noisestate_0/timecount_1[6]  (.D(
        \noisestate_0/timecount_5[6] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[6] ));
    AO1 \state_1ms_0/timecount_RNO_2[3]  (.A(
        \state_1ms_0/PLUSECYCLE[3]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[3] ), 
        .Y(\state_1ms_0/timecount_8_iv_1[3] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[29]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[29]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_482 ));
    DFN1E1 \top_code_0/scaledatain_0[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain_0[0] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_52  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[28] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[10] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[12] ), .Y(
        \timer_top_0/timer_0/N_5 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[14]  (.D(
        \ClockManagement_0/long_timer_0/count_n14 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[14]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m161  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_160 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_161 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_162 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[9] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNI9RKR[1]  (.A(
        \ClockManagement_0/long_timer_0/count[1]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[0]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c1 ));
    XNOR3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m11  (
        .A(\top_code_0_n_divnum_0[2] ), .B(\top_code_0_n_divnum_0[7] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i2_mux ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_12_i ));
    NOR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[3]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_237 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_236 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[3] ));
    OA1B \state_1ms_0/CS_RNO[7]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[7] ), 
        .Y(\state_1ms_0/CS_RNO_3[7] ));
    DFN1E1 \top_code_0/n_divnum[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[9] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_42  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_42_Y ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BFF1_2_inst  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_2_net ));
    AOI1B \DUMP_ON_0/off_on_state_0/state_over_RNO_0  (.A(
        \DUMP_ON_0/off_on_state_0/N_42_i ), .B(
        \DUMP_ON_0/off_on_state_0_state_over ), .C(\DUMP_ON_0/i_5[0] ), 
        .Y(\DUMP_ON_0/off_on_state_0/N_12_mux ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[27]  (.D(
        \top_code_0_dds_configdata[10] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[27]_net_1 ));
    DFN1E1 \top_code_0/scaledatain[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[12] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i18_mux ));
    DFN1 \timer_top_0/state_switch_0/dataout[1]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[1]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[1] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[24]  (.A(
        \DDS_0/dds_state_0/N_305 ), .B(\DDS_0/dds_state_0/N_304 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[24] ), .Y(
        \DDS_0/dds_state_0/N_23 ));
    OR2 OR2_2 (.A(nsctrl_choice_0_dumponoff_rst), .B(net_40), .Y(
        OR2_2_Y));
    DFN1E1 \top_code_0/scaledatain[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[8] ));
    AOI1 \DUMP_OFF_0/off_on_state_0/cs_RNIUSMR[1]  (.A(
        DUMP_OFF_0_dump_off), .B(\DUMP_OFF_0/i_3[1] ), .C(
        \DUMP_OFF_0/off_on_state_0/cs[1]_net_1 ), .Y(
        \DUMP_OFF_0/off_on_state_0/N_42_i ));
    NOR3B \DUMP_0/off_on_state_1/cs_RNO[1]  (.A(
        state1ms_choice_0_reset_out), .B(\DUMP_0/i_0[0] ), .C(
        \DUMP_0/off_on_state_1/N_10 ), .Y(
        \DUMP_0/off_on_state_1/cs_nsss[1] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        );
    MX2C \scalestate_0/CS_RNO_0[2]  (.A(\scalestate_0/CS[2]_net_1 ), 
        .B(\scalestate_0/N_1201 ), .S(timer_top_0_clk_en_scale), .Y(
        \scalestate_0/CS_srsts_i_0[2] ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[10]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[10] ));
    MX2 \noisestate_0/timecount_1_RNO_0[13]  (.A(
        \noisestate_0/acqtime[13]_net_1 ), .B(
        \noisestate_0/dectime[13]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_70 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m22  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_21 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_22 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_23 ));
    NOR2 \scalestate_0/s_acq_RNO_2  (.A(\scalestate_0/CS[4]_net_1 ), 
        .B(\scalestate_0/CS[15]_net_1 ), .Y(
        \scalestate_0/un1_CS6_17_i_a3_0 ));
    DFN1 \timer_top_0/state_switch_0/dataout[10]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[10]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[10] ));
    OR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIQ1684[2]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_2 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE ));
    NOR2B \scalestate_0/timecount_ret_63_RNO_0  (.A(
        \scalestate_0/CUTTIME180[13]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[13] ));
    NOR2B \scalestate_0/CS_RNO[15]  (.A(\scalestate_0/N_1228 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[15]_net_1 ));
    DFN1E1 \top_code_0/pd_pluse_data[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[1] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIARN82[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c6 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c8 ));
    OA1A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_10  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_6 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_7 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_11 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[26]  (.A(
        \DDS_0/dds_state_0/N_472 ), .B(\DDS_0/dds_state_0/N_471 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[26] ), .Y(
        \DDS_0/dds_state_0/N_125 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[8]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[8] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_1[8] ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_12[3]  (.A(
        \DUMP_0/dump_coder_0/para1[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_8[0] ));
    IOPAD_TRI \k2_pad/U0/U0  (.D(\k2_pad/U0/NET1 ), .E(
        \k2_pad/U0/NET2 ), .PAD(k2));
    OA1 \DUMP_0/dump_state_0/cs_RNO[3]  (.A(
        \DUMP_0/dump_state_0/N_196 ), .B(\DUMP_0/dump_state_0/N_195 ), 
        .C(\DUMP_0/dump_state_0/cs4 ), .Y(
        \DUMP_0/dump_state_0/cs_nsss[3] ));
    MX2 \state_1ms_0/timecount_RNO_0[3]  (.A(
        \state_1ms_0/timecount_8[3] ), .B(\state_1ms_0_timecount[3] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_70 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_117  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_117_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[2]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[2]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_487 ));
    MX2 \top_code_0/pluse_str_RNO_0  (.A(top_code_0_pluse_str), .B(
        \top_code_0/un1_xa_49 ), .S(\top_code_0/N_116 ), .Y(
        \top_code_0/N_798 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[0]  (.D(
        \top_code_0_n_divnum_0[0] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[0]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[13]_net_1 ));
    NOR2B \syn_md_module_1/syn_md_0/count_n3_i_a2_0_1  (.A(
        \syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en ), .B(
        top_code_0_scale_rst_3), .Y(\syn_md_module_1/syn_md_0/N_23_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m116  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[19] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_117 ));
    DFN1 \DUMP_0/off_on_timer_0/count[4]  (.D(
        \DUMP_0/off_on_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_2[4] ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_43  (.A(
        \timer_top_0/timer_0/N_8 ), .B(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .Y(
        \timer_top_0/timer_0/I_43 ));
    DFN1E1 \scalestate_0/PLUSETIME180[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[6]_net_1 ));
    NOR2A \plusestate_0/timecount_1_RNO[12]  (.A(\plusestate_0/N_83 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[12] ));
    NOR3A \state_1ms_0/dump_start_RNO_1  (.A(
        \state_1ms_0/un1_CS_9_0_a4_0 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .C(\state_1ms_0/CS[1]_net_1 ), .Y(\state_1ms_0/N_256 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[8] ));
    DFN1 \plusestate_0/dds_config  (.D(
        \plusestate_0/dds_config_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        plusestate_0_dds_config));
    MX2B \PLUSE_0/bri_state_0/cs_RNO[6]  (.A(
        \PLUSE_0/bri_state_0/cs_i_0[6] ), .B(
        \PLUSE_0/bri_state_0/cs[5]_net_1 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_1[6] ));
    DFN1 \top_code_0/relay_on[4]  (.D(
        \top_code_0/relay_on_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[4] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_109  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_133_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_85_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_109_Y ));
    MX2 \noisestate_0/timecount_1_RNO_0[0]  (.A(
        \noisestate_0/acqtime[0]_net_1 ), .B(
        \noisestate_0/dectime[0]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_57 ));
    DFN1 \scalestate_0/rt_sw  (.D(\scalestate_0/rt_sw_RNO_1_net_1 ), 
        .CLK(GLA_net_1), .Q(scalestate_0_rt_sw));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[13]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[13] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[13] ));
    MX2 \scanstate_0/sw_acq2_RNO_0  (.A(scanstate_0_sw_acq2), .B(
        \scanstate_0/N_238 ), .S(\scanstate_0/N_253 ), .Y(
        \scanstate_0/N_109 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[11]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[11] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[11]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i8_mux ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_12_inst  
        (.A(\pd_pluse_top_0/count_0[9] ), .B(
        \pd_pluse_top_0/count_0[10] ), .C(\pd_pluse_top_0/count_0[11] )
        , .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net ));
    NOR2A \DDS_0/dds_state_0/cs_RNO[3]  (.A(\DDS_0/dds_state_0/N_223 ), 
        .B(\DDS_0/dds_state_0/N_227 ), .Y(
        \DDS_0/dds_state_0/cs_RNO[3]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_63_RNO_1  (.A(
        \scalestate_0/OPENTIME[13]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[13] ));
    AO1C \DUMP_0/dump_state_0/cs_i_0_RNI4GHM[0]  (.A(\DUMP_0/i_2[1] ), 
        .B(\DUMP_0/dump_state_0/cs[1]_net_1 ), .C(
        \DUMP_0/dump_state_0/cs_i_0[0]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_171 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/acq_clk  (.A(
        \Signal_Noise_Acq_0/signal_acq_0_Signal_acq_clk ), .B(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .S(
        top_code_0_n_s_ctrl_0), .Y(Signal_Noise_Acq_0_acq_clk));
    AO1 \scalestate_0/timecount_RNO_0[21]  (.A(
        \scalestate_0/CUTTIME180_TEL[21]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[21] )
        , .Y(\scalestate_0/timecount_20_0_iv_0[21] ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[5]_net_1 ));
    NOR2A \scalestate_0/timecount_ret_64_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[13]_net_1 ), .B(\scalestate_0/N_1089 )
        , .Y(\scalestate_0/S_DUMPTIME_m[13] ));
    AX1C 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_2_1_inst  
        (.A(\pd_pluse_top_0/count_6[0] ), .B(
        \pd_pluse_top_0/count_6[1] ), .C(\pd_pluse_top_0/count_6[2] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/count1[2] ));
    MX2 \scanstate_0/timecount_1_RNO_0[13]  (.A(
        \scanstate_0/acqtime[13]_net_1 ), .B(
        \scanstate_0/dectime[13]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_71 ));
    AO1 \PLUSE_0/bri_state_0/cs_RNO_0[1]  (.A(
        \PLUSE_0/bri_state_0/cs[0]_net_1 ), .B(\PLUSE_0/i_3[3] ), .C(
        \PLUSE_0/bri_state_0/cs[2]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/csse_0_0_0_tz ));
    DFN1 \DUMP_0/off_on_state_1/cs[0]  (.D(
        \DUMP_0/off_on_state_1/N_36_i ), .CLK(GLA_net_1), .Q(
        DUMP_0_dump_on));
    DFN1C0 \bridge_div_0/count[1]  (.D(\bridge_div_0/count_5[1] ), 
        .CLK(ddsclkout_c), .CLR(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[1]_net_1 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[1]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_5_2 ), .Y(
        \timer_top_0/timer_0/timedata_4[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m225  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_224 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_225 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_226 ));
    MX2 \scalestate_0/strippluse_RNO_0[6]  (.A(
        \scalestate_0/strippluse_6[6] ), .B(
        \scalestate_0_strippluse[6] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_565 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI1GJG3[12]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c10 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c12 ));
    XA1C \ClockManagement_0/long_timer_0/timeup_RNO_5  (.A(
        \ClockManagement_0/long_timer_0/count[4]_net_1 ), .B(
        \top_code_0_sigtimedata[4] ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_5 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_7 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[19]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[19]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m41_1 ));
    XA1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_7  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[4] )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] )
        );
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/PAND2_20_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc1_25_net ), 
        .C(\sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_17_net ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[15]  (.A(
        \ClockManagement_0/long_timer_0/count_31_0 ), .B(
        \ClockManagement_0/long_timer_0/count[15]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n15 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i6_mux ));
    NOR3B \scanstate_0/CS_i_0_RNI3F711[0]  (.A(\scanstate_0/CS_li[0] ), 
        .B(net_33_0), .C(\scanstate_0/CS[5]_net_1 ), .Y(
        \scanstate_0/timecount_cnst[4] ));
    DFN1E1 \state_1ms_0/CUTTIME[12]  (.D(
        \top_code_0_state_1ms_data[12] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[12]_net_1 ));
    NOR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[8]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_221 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_222 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[8] ));
    NOR2A \timer_top_0/state_switch_0/state_over_n_RNO_3  (.A(
        \timer_top_0/state_switch_0/N_168 ), .B(
        scalestate_0_tetw_pluse), .Y(
        \timer_top_0/state_switch_0/N_280 ));
    DFN1 \DUMP_0/off_on_state_1/cs[1]  (.D(
        \DUMP_0/off_on_state_1/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/off_on_state_1/cs[1]_net_1 ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_3  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_21_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_11_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_17_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_3_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIEP6B[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_9[0] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n15 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI36ES[15]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[15]_net_1 ), .B(
        \sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_15[0] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[4]  (.A(
        \timer_top_0/state_switch_0/N_222 ), .B(
        \timer_top_0/state_switch_0/N_224 ), .C(
        \timer_top_0/state_switch_0/N_223 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[4] ));
    DFN1E1 \scanstate_0/dectime[15]  (.D(\top_code_0_scandata[15] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[15]_net_1 ));
    DFN1 \n_acq_change_0/n_rst_n_0_0  (.D(
        \n_acq_change_0/n_rst_n_0_net_1 ), .CLK(GLA_net_1), .Q(
        n_acq_change_0_n_rst_n_0));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1  (.A(\ADC_c[11] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ));
    XO1 \scalestate_0/M_pulse_RNO_7  (.A(
        \scalestate_0/necount[3]_net_1 ), .B(
        \scalestate_0/M_NUM[3]_net_1 ), .C(\scalestate_0/M_pulse8_1 ), 
        .Y(\scalestate_0/M_pulse8_NE_2 ));
    NOR2B \scalestate_0/load_out_RNO_2  (.A(\scalestate_0/N_1266 ), .B(
        \scalestate_0/N_1251_1 ), .Y(\scalestate_0/un1_CS6_25_i_a3_0 ));
    DFN1E1 \scanstate_0/acqtime[13]  (.D(\top_code_0_scandata[13] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[13]_net_1 ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/i_RNO[4]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[4] ));
    NOR2B \state_1ms_0/timecount_RNO_3[15]  (.A(
        \state_1ms_0/CUTTIME[15]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[15] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n10 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10]/Y ));
    NOR2B \scalestate_0/M_pulse_RNIHCSD  (.A(
        \scalestate_0/timecount_17_sqmuxa_1 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/N_263 ));
    IOPAD_IN \xa_pad[18]/U0/U0  (.PAD(xa[18]), .Y(\xa_pad[18]/U0/NET1 )
        );
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_43  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[3] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[6] ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[10] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        );
    NOR2B \scalestate_0/CS_RNO[6]  (.A(\scalestate_0/N_1221 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO_1[6] ));
    NOR2A \top_code_0/n_s_ctrl_3_i_a2_0  (.A(
        \top_code_0/s_acqnum_1_sqmuxa_1 ), .B(\top_code_0/N_171 ), .Y(
        \top_code_0/N_284 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[11]  (.A(
        \DDS_0/dds_state_0/para[11]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_325 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[11] ));
    DFN1 \scalestate_0/CS[15]  (.D(\scalestate_0/CS_RNO[15]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[15]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[0]  (.A(
        \noisestate_0_timecount[0] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_240 ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_27  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[1] ));
    MX2 \scalestate_0/pn_out_RNO_0  (.A(\scalestate_0/pn_out_4 ), .B(
        scalestate_0_pn_out), .S(\scalestate_0/N_1191 ), .Y(
        \scalestate_0/N_571 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m44_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[15] ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[8]  (.A(
        \top_code_0_dumpdata_0[8] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[8]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[3]  (.A(
        \scalestate_0_timecount[3] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_228 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[6]  (.D(
        \DUMP_0/dump_coder_0/para2_4[6]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[6]_net_1 ));
    IOPAD_BI \xd_pad[11]/U0/U0  (.D(\xd_pad[11]/U0/NET1 ), .E(
        \xd_pad[11]/U0/NET2 ), .Y(\xd_pad[11]/U0/NET3 ), .PAD(xd[11]));
    NOR3B \state_1ms_0/CUTTIME_145_e  (.A(\state_1ms_0/N_16 ), .B(
        \state_1ms_0/un1_PLUSECYCLE13_i_a2_0_net_1 ), .C(
        \top_code_0_state_1ms_lc[0] ), .Y(\state_1ms_0/N_364 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[1]  (.A(\DDS_0/dds_state_0/N_281 )
        , .B(\DDS_0/dds_state_0/N_280 ), .C(
        \DDS_0/dds_state_0/para_9_i_0_1[1] ), .Y(
        \DDS_0/dds_state_0/N_46 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_58  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[28] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[13] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[14] ), .Y(
        \timer_top_0/timer_0/N_3 ));
    DFN1 \state_1ms_0/CS[1]  (.D(\state_1ms_0/CS_RNO_3[1] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[1]_net_1 ));
    AND2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[2] )
        );
    DFN1E1 \DDS_0/dds_state_0/para_reg[6]  (.D(
        \top_code_0_dds_configdata[5] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[6]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[9]  (.D(\GPMI_0_dataout[9] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[9] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_39_i ));
    OA1B \state_1ms_0/CS_RNO[6]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[6] ), 
        .Y(\state_1ms_0/CS_RNO_3[6] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[10] ));
    DFN1E1 \scalestate_0/CUTTIME180[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[9]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[25]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[25]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_309 ));
    NOR2A \PLUSE_0/qq_state_1/Q1Q8_Q2Q7_RNO  (.A(
        \PLUSE_0/qq_state_1/cs4 ), .B(
        \PLUSE_0/qq_state_1/stateover_0_sqmuxa_i_0 ), .Y(
        \PLUSE_0/qq_state_1/Q1Q8_Q2Q7_RNO_0_net_1 ));
    NOR2B \n_acq_change_0/n_acq_start_RNO  (.A(
        \n_acq_change_0/n_acq_start_5 ), .B(net_27), .Y(
        \n_acq_change_0/n_acq_start_RNO_net_1 ));
    DFN1E1 \top_code_0/plusedata[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[3] ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m42_3 ));
    MX2 \scalestate_0/strippluse_RNO_2[9]  (.A(
        \scalestate_0/STRIPNUM180_NUM[9]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[9]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_429 ));
    OR3A \top_code_0/pd_pluse_load_RNO_0  (.A(\xa_c[1] ), .B(
        \top_code_0/N_150 ), .C(\top_code_0/N_167 ), .Y(
        \top_code_0/N_203 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[8]  (.A(
        \plusestate_0_timecount[8] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_249 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[1]  (.A(
        \top_code_0_dumpdata_0[1] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[1] ));
    AOI1B \PLUSE_0/qq_state_1/cs_RNO[1]  (.A(
        \PLUSE_0/qq_state_1/cs_i[0]_net_1 ), .B(
        \PLUSE_0/qq_state_1/N_82 ), .C(\PLUSE_0/qq_state_1/cs4 ), .Y(
        \PLUSE_0/qq_state_1/cs_RNO_2[1] ));
    AND3B 
        \DSTimer_0/dump_sustain_timer_0/cmp_constant_4b_0/AND3B_Temp_0_inst  
        (.A(\DSTimer_0/dump_sustain_timer_0/count[2]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[1]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/cmp_constant_4b_0/Temp_0_net ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[29]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[29]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_483 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[15]  (.A(
        \scanstate_0_timecount[15] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_186 ));
    MX2 \noisestate_0/timecount_1_RNO_0[15]  (.A(
        \noisestate_0/acqtime[15]_net_1 ), .B(
        \noisestate_0/dectime[15]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_72 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m169  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_170 ));
    NOR2B \scalestate_0/timecount_ret_50_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[17]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[17] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[4]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n4 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ));
    MX2 \n_acq_change_0/n_acq_start_RNO_0  (.A(plusestate_0_pluse_acq), 
        .B(noisestate_0_n_acq), .S(top_code_0_pluse_noise_ctrl), .Y(
        \n_acq_change_0/n_acq_start_5 ));
    DFN1E1 \top_code_0/scandata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[7] ));
    DFN1 \ClockManagement_0/clk_10k_0/count[3]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[3] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[3]_net_1 ));
    DFN1E1 \scanstate_0/acqtime[6]  (.D(\top_code_0_scandata[6] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[6]_net_1 ));
    AND3 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_1_8_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_8_net ), 
        .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_8_net ));
    AOI1B \DUMP_0/off_on_state_0/state_over_RNO_0  (.A(
        \DUMP_0/off_on_state_0/N_42_i ), .B(
        \DUMP_0/off_on_state_0_state_over ), .C(\DUMP_0/i_1[0] ), .Y(
        \DUMP_0/off_on_state_0/N_12_mux ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n8 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        );
    MX2 \scalestate_0/strippluse_RNO_0[7]  (.A(
        \scalestate_0/strippluse_6[7] ), .B(
        \scalestate_0_strippluse[7] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_566 ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_3[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_8[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_7[10] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_16[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_19[10] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[1]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[3]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[4]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_492 ));
    OA1B \state_1ms_0/CS_RNO[2]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[2]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[2] ), 
        .Y(\state_1ms_0/CS_RNO_3[2] ));
    NOR3A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_12[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_4[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_7[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_10[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_10[4] ));
    OR2A \plusestate_0/timecount_1_RNO_1[6]  (.A(top_code_0_pluse_rst), 
        .B(\plusestate_0/N_303 ), .Y(\plusestate_0/N_223 ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/i_0[1]  (.A(net_51), .B(net_27)
        , .Y(\i_0_0[1] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[1]  (.A(
        \DDS_0/dds_state_0/para[1]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569 ), .C(\DDS_0/dds_state_0/N_278 ), .Y(
        \DDS_0/dds_state_0/para_9_i_0_1[1] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m46_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[13] ));
    AND3 \scalestate_0/necount_inc_0/AND2_6_inst  (.A(
        \scalestate_0/necount[3]_net_1 ), .B(
        \scalestate_0/necount[4]_net_1 ), .C(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/inc_5_net ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[0]  (.D(
        \top_code_0_bri_datain[4] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[0] ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_12  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_3 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[13]  (.A(
        \plusestate_0_timecount[13] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_194 ));
    MX2 \scalestate_0/strippluse_RNO_2[0]  (.A(
        \scalestate_0/STRIPNUM180_NUM[0]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[0]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_420 ));
    OA1B \PLUSE_0/bri_state_0/up_RNO_0  (.A(
        \PLUSE_0/bri_state_0/cs[1]_net_1 ), .B(
        \PLUSE_0/bri_state_0/N_179 ), .C(\PLUSE_0/i_3[2] ), .Y(
        \PLUSE_0/bri_state_0/N_178 ));
    AO1A \scalestate_0/timecount_ret_37_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[3]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[3] ), .Y(
        \scalestate_0/timecount_20_iv_1[3] ));
    DFN1 \top_code_0/state_1ms_start_ret_3  (.D(\top_code_0/N_112 ), 
        .CLK(GLA_net_1), .Q(\top_code_0/N_112_reto ));
    OR3A \scalestate_0/reset_out_RNO_1  (.A(\scalestate_0/N_1208 ), .B(
        \scalestate_0/CS_0[11]_net_1 ), .C(
        \scalestate_0/un1_CS_44_i_0 ), .Y(\scalestate_0/N_1097 ));
    DFN1 \plusestate_0/CS[9]  (.D(\plusestate_0/CS_RNO[9]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[9]_net_1 ));
    DFN1E0 \DDS_0/dds_state_0/para[7]  (.D(\DDS_0/dds_state_0/N_8 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[7]_net_1 ));
    DFN1E1 \scanstate_0/timecount_1[15]  (.D(
        \scanstate_0/timecount_5[15] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[15] ));
    NOR2A \top_code_0/n_divnum_1_sqmuxa_0_a2_0  (.A(\top_code_0/N_329 )
        , .B(\top_code_0/N_150 ), .Y(\top_code_0/N_339 ));
    MX2A \scalestate_0/off_test_RNO_0  (.A(\scalestate_0/N_1262 ), .B(
        scalestate_0_off_test), .S(\scalestate_0/N_1175 ), .Y(
        \scalestate_0/N_726 ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[5]  (.A(
        \PLUSE_0/bri_state_0/cs[5]_net_1 ), .B(
        \PLUSE_0/bri_state_0/csse_4_0_a4_0_0 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[5] ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i2_mux ));
    OR2A \top_code_0/s_acqnum_1_sqmuxa_0_o2_0  (.A(\xa_c[2] ), .B(
        \xa_c[3] ), .Y(\top_code_0/N_142 ));
    NOR2B \top_code_0/relay_on_RNO[6]  (.A(\top_code_0/N_815 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[6]_net_1 ));
    NOR3B \top_code_0/dump_cho_1_sqmuxa_0_a2  (.A(\top_code_0/N_331 ), 
        .B(\top_code_0/N_334 ), .C(\top_code_0/N_147 ), .Y(
        \top_code_0/dump_cho_1_sqmuxa ));
    AO1 \state_1ms_0/timecount_RNO_4[4]  (.A(
        \state_1ms_0/S_DUMPTIME[4]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[4] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[4] ));
    NOR3C \DUMP_ON_0/off_on_coder_0/i_RNO[1]  (.A(
        \DUMP_ON_0/off_on_coder_0/i_0_2[1] ), .B(
        \DUMP_ON_0/off_on_coder_0/i_0_1[1] ), .C(OR2_2_Y), .Y(
        \DUMP_ON_0/off_on_coder_0/i_RNO_5[1] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[3]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n3 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ));
    IOPAD_IN \gpio_pad/U0/U0  (.PAD(gpio), .Y(\gpio_pad/U0/NET1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[5]  (.A(
        \s_acq_change_0/s_stripnum_5[5] ), .B(
        \s_acq_change_0_s_stripnum[5] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_61 ));
    DFN1E1 \top_code_0/cal_data[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[3] ));
    CLKINT \s_acq_change_0/s_rst_RNIKACF  (.A(
        \s_acq_change_0/s_rst_net_1 ), .Y(s_acq_change_0_s_rst));
    AO1A \plusestate_0/off_test_RNO_0  (.A(\plusestate_0/CS[5]_net_1 ), 
        .B(plusestate_0_off_test), .C(\plusestate_0/CS[4]_net_1 ), .Y(
        \plusestate_0/N_141 ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ));
    DFN1E1 \scalestate_0/DUMPTIME[2]  (.D(\top_code_0_scaledatain[2] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[2]_net_1 ));
    DFN1E0 \DDS_0/dds_state_0/para[12]  (.D(\DDS_0/dds_state_0/N_103 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[12]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[7]  (.D(\top_code_0_scaledatain[7] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[7]_net_1 ));
    NOR2A \DUMP_0/off_on_timer_0/count_RNO[0]  (.A(
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_0/count_2[0] ), .Y(\DUMP_0/off_on_timer_0/count_n0 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[2] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[12]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[12] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count[12] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[0]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[0] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_6[0] ));
    NOR2A \noisestate_0/timecount_1_RNO[1]  (.A(\noisestate_0/N_58 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[1] ));
    NOR3A \timer_top_0/state_switch_0/state_start5_0_0_a2_0_1  (.A(
        top_code_0_scale_start), .B(top_code_0_scan_start), .C(
        top_code_0_noise_start), .Y(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_0_0 ));
    NOR2B \scalestate_0/timecount_ret_11_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[7]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[7] ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[10]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[10] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_10_inst ), .S(top_code_0_n_s_ctrl_0)
        , .Y(\Signal_Noise_Acq_0_dataout[10] ));
    OR3 \scalestate_0/timecount_ret_67_RNO  (.A(
        \scalestate_0/ACQTIME_m[14] ), .B(
        \scalestate_0/PLUSETIME90_m[14] ), .C(
        \scalestate_0/S_DUMPTIME_m[14] ), .Y(
        \scalestate_0/timecount_20_iv_6[14] ));
    DFN1 \plusestate_0/CS[5]  (.D(\plusestate_0/CS_RNO_0[5]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[5]_net_1 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_14  (.A(\xd_in[0] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[0] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n11 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        );
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNI18A22[6]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c4 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c6 ));
    NOR2 \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[10]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 ), .B(
        \pd_pluse_top_0/i_1[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_180 ));
    DFN1E1 \top_code_0/dump_cho[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/dump_cho_1_sqmuxa ), .Q(
        \top_code_0_dump_cho_0[1] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_31  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_31_Y ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI8SKV[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_5[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_7[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_3[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_9[0] ));
    NOR2 \pd_pluse_top_0/pd_pluse_state_0/cs_RNIFFJJ[4]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[4]_net_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[7]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_srsts_0_i_a5_1[12] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[12]  (.A(
        \scanstate_0_timecount[12] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_256 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[0]_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[22]  (.D(
        \top_code_0_dds_configdata[5] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[22]_net_1 ));
    NOR3B \timer_top_0/state_switch_0/state_start5_0_0_a2_2  (.A(
        \timer_top_0/state_switch_0/N_284 ), .B(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_2_0_net_1 ), 
        .C(top_code_0_scale_start), .Y(
        \timer_top_0/state_switch_0/N_296 ));
    DFN1 \timer_top_0/state_switch_0/state_over_n  (.D(
        \timer_top_0/state_switch_0/N_78 ), .CLK(GLA_net_1), .Q(
        \timer_top_0/state_switch_0_state_over_n ));
    AO1 \scalestate_0/timecount_ret_11_RNO_2  (.A(
        \scalestate_0/CUTTIME180[7]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[7] ), .Y(
        \scalestate_0/timecount_20_iv_2[7] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[13]  (.A(
        \DDS_0/dds_state_0/para[13]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_334 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[13] ));
    OR2B \DUMP_OFF_1/off_on_state_0/state_over_RNO  (.A(
        \DUMP_OFF_1/off_on_state_0/N_12_mux ), .B(
        nsctrl_choice_0_dumponoff_rst), .Y(
        \DUMP_OFF_1/off_on_state_0/N_9 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n4 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4]/Y ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/QXOR2_16_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_20_net ), 
        .B(\sd_acq_top_0/count[20] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[20] ));
    NOR3C \scalestate_0/timecount_ret_85_RNO_0  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[11]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[11] ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[11]  (.D(
        \ClockManagement_0/long_timer_0/count_n11 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[11]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[0] ));
    DFN1E1 \top_code_0/s_acqnum[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[11] ));
    IOPAD_BI \xd_pad[12]/U0/U0  (.D(\xd_pad[12]/U0/NET1 ), .E(
        \xd_pad[12]/U0/NET2 ), .Y(\xd_pad[12]/U0/NET3 ), .PAD(xd[12]));
    DFN1 \DSTimer_0/dump_sustain_timer_0/data[0]  (.D(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[0]_net_1 ), .CLK(
        GLA_net_1), .Q(\DSTimer_0/dump_sustain_timer_0/data[0]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[8]_net_1 ));
    DFN1 \scalestate_0/s_acqnum_1[8]  (.D(
        \scalestate_0/s_acqnum_1_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[8] ));
    XOR2 \PLUSE_0/bri_timer_0/count_RNO[3]  (.A(
        \PLUSE_0/bri_timer_0/count_c2 ), .B(\PLUSE_0/count_8[3] ), .Y(
        \PLUSE_0/bri_timer_0/count_n3 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[28]  (.A(
        \DDS_0/dds_state_0/N_480 ), .B(\DDS_0/dds_state_0/N_479 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[28] ), .Y(
        \DDS_0/dds_state_0/N_129 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[7]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[2]_net_1 ));
    NOR3B \DUMP_0/off_on_coder_0/i_RNO_0[1]  (.A(\DUMP_0/count_0[4] ), 
        .B(\DUMP_0/count_0[2] ), .C(\DUMP_0/count_0[3] ), .Y(
        \DUMP_0/off_on_coder_0/i_0_2[1] ));
    NOR3C \sd_acq_top_0/sd_sacq_state_0/cs_RNO[11]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[10]_net_1 ), .B(
        \sd_acq_top_0/i_0[8] ), .C(\sd_acq_top_0/sd_sacq_state_0/cs4 ), 
        .Y(\sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[11] ));
    DFN1E1 \top_code_0/state_1ms_data[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[10] ));
    NOR2B \timer_top_0/state_switch_0/clk_en_pluse_RNO  (.A(
        \timer_top_0/state_switch_0/N_293 ), .B(
        \timer_top_0/timer_0_time_up ), .Y(
        \timer_top_0/state_switch_0/clk_en_pluse_RNO_net_1 ));
    XOR2 \PLUSE_0/qq_coder_0/un1_qq_para2_2[0]  (.A(
        \PLUSE_0/qq_para2[2] ), .B(\PLUSE_0/count_9[2] ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_2[0]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_41_i ));
    NOR3C \scalestate_0/timecount_RNO_3[21]  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[21]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[21] ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[9]  (.D(
        \top_code_0_state_1ms_data[9] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[9]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[4]  (.D(\GPMI_0_dataout_0[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[4] ));
    DFN1E1 \top_code_0/scandata[14]  (.D(\GPMI_0_dataout[14] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[14] ));
    OR3 \top_code_0/dds_choice_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_161 ), .Y(
        \top_code_0/N_205 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m87  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_88 ));
    DFN1E1 \scanstate_0/acqtime[14]  (.D(\top_code_0_scandata[14] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[14]_net_1 ));
    DFN1 \top_code_0/noise_start_ret_2  (.D(\top_code_0/un1_xa_13 ), 
        .CLK(GLA_net_1), .Q(\top_code_0/un1_xa_13_reto ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[21]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[21]_net_1 ));
    IOIN_IB \xa_pad[10]/U0/U1  (.YIN(\xa_pad[10]/U0/NET1 ), .Y(
        \xa_c[10] ));
    DFN1E1 \top_code_0/scalechoice[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0[1] ));
    OR3 \state_1ms_0/timecount_RNO_1[7]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[7] ), .B(
        \state_1ms_0/CUTTIME_m[7] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[7] ), .Y(
        \state_1ms_0/timecount_8[7] ));
    DFN1E1 \top_code_0/bri_datain[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[9] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[16]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[16]_net_1 ));
    NOR3C \scalestate_0/timecount_20_iv_5_RNO_1[5]  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[5]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[5] ));
    OR2A \scalestate_0/necount_cmp_0/OR2A_4  (.A(
        \scalestate_0/necount[2]_net_1 ), .B(
        \scalestate_0/M_NUM[2]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_4_Y ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datatwo  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ));
    DFN1 \scalestate_0/necount[6]  (.D(
        \scalestate_0/necount_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[6]_net_1 ));
    DFN1E1 \top_code_0/cal_data[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[1] ));
    NOR2B \noisestate_0/dumpon_ctr_RNO  (.A(\noisestate_0/N_130 ), .B(
        top_code_0_noise_rst), .Y(\noisestate_0/dumpon_ctr_RNO_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[8]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIOH1G[2]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[2]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_2[0] ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/data_RNO[3]  (.A(
        \DSTimer_0/dump_sustain_timer_0/N_27 ), .B(
        top_code_0_dump_sustain), .Y(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[3]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/dataout[15]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[15] ), .B(
        top_code_0_n_s_ctrl_1), .Y(\Signal_Noise_Acq_0_dataout[15] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI7G3A[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_6[0] ));
    IOTRI_ORE_EB \rt_sw_pad/U0/U1  (.D(\state1ms_choice_0/rt_sw_4 ), 
        .E(VCC), .OCE(net_27), .OCLK(GLA_net_1), .DOUT(
        \rt_sw_pad/U0/NET1 ), .EOUT(\rt_sw_pad/U0/NET2 ));
    AO1 \scalestate_0/timecount_20_iv_4[4]  (.A(
        \scalestate_0/CUTTIMEI90[4]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[4] ), .Y(
        \scalestate_0/timecount_20_iv_4[4]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m131  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[19] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_132 ));
    DFN1 \DUMP_0/dump_state_0/cs[3]  (.D(
        \DUMP_0/dump_state_0/cs_nsss[3] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[3]_net_1 ));
    AO1C \state_1ms_0/CS_RNO_0[5]  (.A(\state_1ms_0/CS[4]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[5] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m11  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_8_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_11_0 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_12_0 ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/enable  (.A(
        scalestate_0_dump_sustain_ctrl), .B(top_code_0_dump_sustain), 
        .Y(\DSTimer_0/dump_sustain_timer_0/enable_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI16T7[4]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_4[0] ));
    DFN1C0 \bridge_div_0/count[4]  (.D(\bridge_div_0/count_5[4] ), 
        .CLK(ddsclkout_c), .CLR(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[4]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/ADD_20x20_slow_I19_Y_2 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[19] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_1_8_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_8_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_8_net ));
    NOR2B \scalestate_0/s_acq_RNO  (.A(\scalestate_0/N_724 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/s_acq_RNO_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[6]  (.D(
        \DUMP_0/dump_coder_0/para4_4[6]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[6]_net_1 ));
    DFN1E1 \top_code_0/noisedata[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[10] ));
    DFN1E1 \scalestate_0/CUTTIME90[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_134  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_134_Y ));
    DFN1E1 \plusestate_0/timecount_1[9]  (.D(
        \plusestate_0/timecount_5[9] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[9] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[3]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[3]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_491 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[16]  (.D(
        \top_code_0_dds_configdata[15] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[16]_net_1 ));
    MX2 \scalestate_0/necount_RNO_0[2]  (.A(\scalestate_0/necount1[2] )
        , .B(\scalestate_0/necount[2]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_732 ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIMR3H2[6]  (.A(
        \DUMP_0/dump_timer_0/count_c5 ), .B(\DUMP_0/count_0[6] ), .Y(
        \DUMP_0/dump_timer_0/count_c6 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i22_mux ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_4  (.A(
        \scalestate_0/necount[10]_net_1 ), .B(
        \scalestate_0/M_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_4_Y ));
    NOR2B \ClockManagement_0/clk_10k_0/un1_count_1_I_42  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_1[0] ), 
        .Y(\ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_11[0] ));
    OR2A \top_code_0/un1_state_1ms_rst_n117_4_i_o2  (.A(\xa_c[3] ), .B(
        \xa_c[1] ), .Y(\top_code_0/N_161 ));
    OR2A \noisestate_0/sw_acq2_RNO  (.A(top_code_0_noise_rst), .B(
        \noisestate_0/N_108 ), .Y(\noisestate_0/sw_acq2_RNO_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIEKR21[21]  (.A(
        \sd_acq_top_0/count[21] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[21]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_17[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_0[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[1]_net_1 ));
    NOR2B \bri_dump_sw_0/dump_start_RNO  (.A(
        \bri_dump_sw_0/dump_start_5 ), .B(net_27), .Y(
        \bri_dump_sw_0/dump_start_RNO_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[15]  (.A(
        \scalestate_0_timecount[15] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_188 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[11]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[11]_net_1 ), .CLK(
        ddsclkout_c), .Q(
        \pd_pluse_top_0/pd_pluse_state_0/cs[11]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs_i[0]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .CLK(ddsclkout_c), .Q(
        \sd_acq_top_0/sd_sacq_state_0/cs_i[0]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[9]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[9]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_288 ));
    DFN1E0 \DDS_0/dds_state_0/para[28]  (.D(\DDS_0/dds_state_0/N_129 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[28]_net_1 ));
    AO1 \scalestate_0/timecount_RNO_2[20]  (.A(
        \scalestate_0/CUTTIMEI90[20]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[20] ), .Y(
        \scalestate_0/timecount_20_0_iv_1[20] ));
    DFN1E0 \DDS_0/dds_state_0/para[17]  (.D(\DDS_0/dds_state_0/N_161 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[17]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[19]  (.A(
        \scalestate_0_timecount[19] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_272 ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_5 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_9 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m115  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_114 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_115 ), .S(
        \top_code_0_s_addchoice_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_116 ));
    NOR2B \scanstate_0/acqtime_0_sqmuxa  (.A(top_code_0_scanchoice), 
        .B(top_code_0_scanload), .Y(
        \scanstate_0/acqtime_0_sqmuxa_net_1 ));
    MX2 \state_1ms_0/timecount_RNO_0[14]  (.A(
        \state_1ms_0/timecount_8[14] ), .B(\state_1ms_0_timecount[14] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_81 ));
    NOR3C \scalestate_0/timecount_ret_8_RNO_1  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[3]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[3] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/QAND2_26_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net ), 
        .C(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_31_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_20_net ));
    DFN1E1 \top_code_0/noisedata[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[3] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[10]_net_1 )
        );
    DFN1E0 \DUMP_0/dump_coder_0/para2[10]  (.D(
        \DUMP_0/dump_coder_0/para2_4[10]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[10]_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_66_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 )
        , .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_3_i_a2_1 ), 
        .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_14[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[14]_net_1 ), .B(
        \sd_acq_top_0/count_0[14] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_14[0] ));
    AO1 \syn_md_module_1/syn_md_0/count_RNO_1[2]  (.A(
        \syn_md_module_1/syn_md_0/count_n2_i_a2_0 ), .B(
        top_code_0_scale_rst_2), .C(\syn_md_module_1/syn_md_0/N_23_1 ), 
        .Y(\syn_md_module_1/syn_md_0/count_n2_i_0 ));
    MX2 \scanstate_0/soft_d_RNO_0  (.A(scanstate_0_soft_d), .B(
        \scanstate_0/CS[1]_net_1 ), .S(\scanstate_0/N_253 ), .Y(
        \scanstate_0/N_110 ));
    DFN1E1 \scalestate_0/NE_NUM[1]  (.D(\top_code_0_scaledatain[1] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[1]_net_1 ));
    DFN1E1 \top_code_0/scaledatain[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[6] ));
    DFN1E1 \scalestate_0/CUTTIME90[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[14]_net_1 ));
    NOR3B \top_code_0/relay_close_1_sqmuxa_0_a2  (.A(\xa_c[6] ), .B(
        \top_code_0/relay_close_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_137 ), .Y(\top_code_0/relay_close_1_sqmuxa ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[2]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n2 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ));
    DFN1E1 \top_code_0/state_1ms_load  (.D(\top_code_0/N_106 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_state_1ms_load));
    NOR2 \DUMP_0/off_on_coder_0/i_RNO_1[1]  (.A(\DUMP_0/count_0[1] ), 
        .B(\DUMP_0/count_0[0] ), .Y(\DUMP_0/off_on_coder_0/i_0_1[1] ));
    DFN1E1 \top_code_0/dds_configdata[4]  (.D(\GPMI_0_dataout[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[4] ));
    NOR2B \scalestate_0/timecount_ret_90_RNO_0  (.A(
        \scalestate_0/OPENTIME[8]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[8] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[4]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[2]  (.D(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[2] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/i_1[2] ));
    NOR2B \scanstate_0/dumpoff_ctr_RNO  (.A(\scanstate_0/N_113 ), .B(
        net_33), .Y(\scanstate_0/dumpoff_ctr_RNO_3 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m207  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_206 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_207 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_208 ));
    NOR2B \scalestate_0/timecount_ret_53_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[18]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[18] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_54_i ));
    DFN1E1 \top_code_0/sigtimedata[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[9] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_64_i ));
    NOR3C \scalestate_0/timecount_ret_63_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[13]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[13] ));
    DFN1E1 \scalestate_0/ACQ180_NUM[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[11]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[9]_net_1 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_3_inst  
        (.A(\pd_pluse_top_0/count_6[0] ), .B(
        \pd_pluse_top_0/count_6[1] ), .C(\pd_pluse_top_0/count_6[2] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net ));
    XOR2 \ClockManagement_0/clk_div500_0/un1_count_1_I_33  (.A(
        \ClockManagement_0/clk_div500_0/count[1]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_TMP[0] ), .Y(
        \ClockManagement_0/clk_div500_0/I_33 ));
    MX2 \scalestate_0/strippluse_RNO_2[6]  (.A(
        \scalestate_0/STRIPNUM180_NUM[6]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[6]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_426 ));
    MX2 \top_code_0/relay_on_RNO_0[7]  (.A(\relay_on_c[7] ), .B(
        \GPMI_0_dataout[7] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_816 ));
    NOR2B \state_1ms_0/timecount_RNO_3[9]  (.A(
        \state_1ms_0/CUTTIME[9]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[9] ));
    DFN1E1 \top_code_0/dumpdata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[7] ));
    XA1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_41  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_48_i ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] )
        );
    DFN1E1 \scalestate_0/NE_NUM[7]  (.D(\top_code_0_scaledatain[7] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[7]_net_1 ));
    AO1B \plusestate_0/pluse_acq_RNO_0  (.A(plusestate_0_pluse_acq), 
        .B(\plusestate_0/N_302 ), .C(\plusestate_0/N_305 ), .Y(
        \plusestate_0/N_122 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_6[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[1]_net_1 ), .B(
        \pd_pluse_top_0/count_6[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_1[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m60  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_59 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_60 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_61 ));
    MX2 \state_1ms_0/timecount_RNO_0[12]  (.A(
        \state_1ms_0/timecount_8[12] ), .B(\state_1ms_0_timecount[12] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_79 ));
    IOPAD_TRI \ddsdata_pad/U0/U0  (.D(\ddsdata_pad/U0/NET1 ), .E(
        \ddsdata_pad/U0/NET2 ), .PAD(ddsdata));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[5]  (.D(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[5] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/i_0[5] ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[6]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_34 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[6] ));
    NOR2B \state_1ms_0/timecount_RNO[9]  (.A(\state_1ms_0/N_76 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[9]_net_1 ));
    MX2 \plusestate_0/timecount_1_RNO[3]  (.A(\plusestate_0/N_74 ), .B(
        \plusestate_0/timecount_cnst[3] ), .S(\plusestate_0/N_271 ), 
        .Y(\plusestate_0/timecount_5[3] ));
    DFN1 \top_code_0/relay_on[9]  (.D(
        \top_code_0/relay_on_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[9] ));
    NOR2B \state_1ms_0/timecount_RNO_5[8]  (.A(
        \state_1ms_0/PLUSECYCLE[8]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[8] ));
    NOR2B \nsctrl_choice_0/dumponoff_rst_RNO  (.A(
        \nsctrl_choice_0/dumponoff_rst_5 ), .B(net_27), .Y(
        \nsctrl_choice_0/dumponoff_rst_RNO_net_1 ));
    OA1C \top_code_0/nstateload_RNO  (.A(\top_code_0/N_211 ), .B(
        top_code_0_nstateload), .C(\top_code_0/N_288 ), .Y(
        \top_code_0/N_80 ));
    OR3 \topctrlchange_0/soft_dump_6_iv  (.A(
        \topctrlchange_0/s_dumpin2_m ), .B(
        \topctrlchange_0/s_dumpin3_m ), .C(
        \topctrlchange_0/s_dumpin1_m ), .Y(
        \topctrlchange_0/soft_dump_6 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m190  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_191 ));
    AX1C \scalestate_0/necount_inc_0/XOR2_3_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount[3]_net_1 ), .C(
        \scalestate_0/necount[4]_net_1 ), .Y(
        \scalestate_0/necount1[4] ));
    DFN1E1 \plusestate_0/PLUSETIME[14]  (.D(\top_code_0_plusedata[14] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[14]_net_1 ));
    NOR3 \top_code_0/pd_pluse_load_RNO_1  (.A(\top_code_0/N_150 ), .B(
        \top_code_0/N_167 ), .C(\top_code_0/N_157 ), .Y(
        \top_code_0/N_290 ));
    DFN1E0 \DDS_0/dds_state_0/para[26]  (.D(\DDS_0/dds_state_0/N_125 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[26]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_4_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_4_net ));
    XOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIMN7R[4]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[4]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_4 ));
    DFN1E1 \top_code_0/sd_sacq_data[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[9] ));
    IOPAD_TRI \Q3Q6_pad/U0/U0  (.D(\Q3Q6_pad/U0/NET1 ), .E(
        \Q3Q6_pad/U0/NET2 ), .PAD(Q3Q6));
    DFN1E1 \state_1ms_0/PLUSECYCLE[10]  (.D(
        \top_code_0_state_1ms_data[10] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[10]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_57  (.D(
        \scalestate_0/timecount_20_iv_7[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[0] ));
    AO1C \DUMP_0/dump_coder_0/un1_para114_4  (.A(
        \DUMP_0/dump_coder_0/para17_net_1 ), .B(
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ), .C(
        top_code_0_dumpload), .Y(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[17]  (.D(
        \top_code_0_dds_configdata[0] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[17]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[2]  (.A(
        \state_1ms_0_timecount[2] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_232 ));
    NOR3C \scalestate_0/timecount_ret_53_RNO_1  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[18]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[18] ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_2  (.A(
        \scalestate_0/NE_NUM[8]_net_1 ), .B(
        \scalestate_0/necount[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_2_Y ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[12]  (.A(
        \scalestate_0_timecount[12] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_258 ));
    OR3 \scalestate_0/timecount_ret_73_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[7] ), .B(
        \scalestate_0/OPENTIME_TEL_m[7] ), .C(
        \scalestate_0/timecount_20_iv_4[7] ), .Y(
        \scalestate_0/timecount_20_iv_8[7] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_21[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_4[0] ));
    AO1A \state_1ms_0/timecount_RNO_2[6]  (.A(
        \state_1ms_0/PLUSECYCLE[6]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/PLUSETIME_i_m[6] ), 
        .Y(\state_1ms_0/timecount_8_iv_1[6] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[18]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[18]_net_1 ));
    AX1C \ClockManagement_0/clk_10k_0/un1_count_1_I_32  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \ClockManagement_0/clk_10k_0/count[4]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/I_32_0 ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y ));
    IOPAD_IN \xa_pad[8]/U0/U0  (.PAD(xa[8]), .Y(\xa_pad[8]/U0/NET1 ));
    NOR2A \scalestate_0/CS_RNID9K6[14]  (.A(\scalestate_0/N_1262 ), .B(
        \scalestate_0/CS[14]_net_1 ), .Y(\scalestate_0/N_1266 ));
    NOR3C \ClockManagement_0/clk_10k_0/un1_count_1_I_49  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_1[0] ), 
        .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_2[0] ), 
        .C(\ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] ), 
        .Y(\ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_3[0] ));
    NOR2B \scalestate_0/necount_RNO[8]  (.A(\scalestate_0/N_738 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[8]_net_1 ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_3  (.A(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .B(
        \timer_top_0/dataout[13] ), .C(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_3_Y ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNILOCG[7]  (.A(
        \DUMP_0/dump_coder_0/para2[7]_net_1 ), .B(\DUMP_0/count_0[7] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_7[0] ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[2]  (.A(
        \Signal_Noise_Acq_0/un1_signal_acq_0[2] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_2_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[2] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[5]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[12]_net_1 ));
    DFN1P0 \bridge_div_0/count[0]  (.D(\bridge_div_0/count_5[0] ), 
        .CLK(ddsclkout_c), .PRE(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[0]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_58_i ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[7]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[7] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_3[7] ));
    AO1C \scalestate_0/s_acq_RNO_1  (.A(\scalestate_0/N_1197 ), .B(
        \scalestate_0/un1_CS6_17_i_a3_0 ), .C(
        timer_top_0_clk_en_scale_0), .Y(\scalestate_0/N_1169 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m20  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_21 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[7]  (.A(
        \s_acq_change_0/s_acqnum_5[7] ), .B(
        \s_acq_change_0_s_acqnum[7] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_77 ));
    NOR2B \scalestate_0/M_pulse_RNO  (.A(\scalestate_0/N_745 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/M_pulse_RNO_net_1 ));
    DFN1E1 \top_code_0/noisedata[12]  (.D(\GPMI_0_dataout[12] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[12] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[10]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[10] ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_5  (.A(
        \scalestate_0/necount[5]_net_1 ), .B(
        \scalestate_0/NE_NUM[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_5_Y ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[1]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[1] ));
    DFN1 \top_code_0/relay_close[0]  (.D(
        \top_code_0/relay_close_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[0] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[13]  (.A(
        \s_acq_change_0/s_acqnum_5[13] ), .B(
        \s_acq_change_0_s_acqnum[13] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_83 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m139  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[3] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_140 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_2_i ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[24]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[24]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_303 ));
    XA1A \ClockManagement_0/long_timer_0/timeup_RNO_4  (.A(
        \ClockManagement_0/long_timer_0/count[15]_net_1 ), .B(
        \top_code_0_sigtimedata[15] ), .C(
        \ClockManagement_0/long_timer_0/clk_5K_en_1 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_0 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2b_12_inst  (
        .A(\sd_acq_top_0/count_10[3] ), .B(\sd_acq_top_0/count_10[4] ), 
        .C(\sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_5_net ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m151  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_152 ));
    OR3 \DUMP_0/dump_coder_0/para6_RNI4RMA8[0]  (.A(
        \DUMP_0/dump_coder_0/i_reg16_NE_7[0] ), .B(
        \DUMP_0/dump_coder_0/i_reg16_NE_6[0] ), .C(
        \DUMP_0/dump_coder_0/i_reg16_NE_8[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE[0] ));
    AO1A \scalestate_0/timecount_ret_77_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[6]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[6] ), .Y(
        \scalestate_0/timecount_20_iv_0[6] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIRIUE[4]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[4]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_4[0] ));
    NOR2A \scanstate_0/timecount_1_RNO[14]  (.A(\scanstate_0/N_72 ), 
        .B(\scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[14] ));
    DFN1E1 \bridge_div_0/datahalf[0]  (.D(\top_code_0_scaleddsdiv[0] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/datahalf[0]_net_1 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[0]  (.A(\s_acq_change_0/N_56 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[0]_net_1 ));
    NOR2A \timer_top_0/timer_0/Timer_Cmp_0/NOR2A_0  (.A(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .B(
        \timer_top_0/dataout[20] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR2A_0_Y ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_11_0  (.A(\xd_in[3] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout_0[3] ));
    DFN1 \noisestate_0/n_acq  (.D(\noisestate_0/n_acq_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(noisestate_0_n_acq));
    DFN1 \timer_top_0/state_switch_0/dataout[14]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[14]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[14] ));
    DFN1E1 \scalestate_0/PLUSETIME180[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[11]_net_1 ));
    NOR2A \plusestate_0/timecount_1_RNO[9]  (.A(\plusestate_0/N_80 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[9] ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[6]_net_1 ));
    DFN1 \n_acq_change_0/n_rst_n  (.D(\n_acq_change_0/n_rst_n_0_net_1 )
        , .CLK(GLA_net_1), .Q(n_acq_change_0_n_rst_n));
    DFN1 \top_code_0/dump_sustain  (.D(
        \top_code_0/dump_sustain_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        top_code_0_dump_sustain));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_50_i ));
    IOPAD_BI \xd_pad[14]/U0/U0  (.D(\xd_pad[14]/U0/NET1 ), .E(
        \xd_pad[14]/U0/NET2 ), .Y(\xd_pad[14]/U0/NET3 ), .PAD(xd[14]));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para1[1]  (.D(
        \top_code_0_bri_datain[1] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para1[1] ));
    NOR2B \scalestate_0/timecount_20_iv_5_RNO_0[11]  (.A(
        \scalestate_0/OPENTIME_TEL[11]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[11] ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_31  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_42_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[7] )
        );
    DFN1E1 \scalestate_0/ACQECHO_NUM[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[9]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m287  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_288 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[3]  (.D(
        \top_code_0_dds_configdata[2] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[3]_net_1 ));
    DFN1E1 \noisestate_0/dectime[7]  (.D(\top_code_0_noisedata[7] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[7]_net_1 ));
    XOR2 \ClockManagement_0/clk_div500_0/un1_count_1_I_23  (.A(
        \ClockManagement_0/clk_div500_0/count[0]_net_1 ), .B(
        \ClockManagement_0/clk_5M_en ), .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_partial_sum[0] )
        );
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I7_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I6_un1_CO1 ), 
        .B(\s_acq_change_0_s_stripnum[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N160 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m84  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_85 ));
    DFN1E1 \top_code_0/scaleddsdiv[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[5] ));
    DFN1E1 \top_code_0/pd_pluse_data[6]  (.D(\GPMI_0_dataout[6] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[6] ));
    NOR3C \scalestate_0/timecount_ret_28_RNO_3  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[1]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[1] ));
    DFN1E1 \top_code_0/scandata[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[0] ));
    DFN1E1 \scalestate_0/timecount_ret_52  (.D(
        \scalestate_0/OPENTIME_TEL_m[18] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/OPENTIME_TEL_m_reto[18] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[4]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[4] ));
    DFN1E1 \top_code_0/sigtimedata[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[2] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m68  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_69 ));
    NOR2B \scalestate_0/timecount_ret_71_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[15]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[15] ));
    DFN1E1 \noisestate_0/timecount_1[8]  (.D(
        \noisestate_0/timecount_5[8] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[8] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_157  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_24_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_121_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_157_Y ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIOUJ12[2]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_12[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_2[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_5[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_10[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m205  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[9] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_206 ));
    NOR2B \scalestate_0/timecount_ret_28_RNO_4  (.A(
        \scalestate_0/OPENTIME[1]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[1] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[12]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[11] )
        , .Y(\DDS_0/dds_state_0/N_329 ));
    DFN1E1 \top_code_0/sigtimedata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[7] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[2] ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_1  (.A(
        \scalestate_0/NE_NUM[10]_net_1 ), .B(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_1_Y ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[10]  (.A(
        \scalestate_0/s_acqnum_7[10] ), .B(\scalestate_0_s_acqnum[10] )
        , .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_557 ));
    NOR2B \scalestate_0/necount_LE_M_RNINMTM  (.A(
        \scalestate_0/timecount_13_sqmuxa_0 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/N_259 ));
    DFN1 \DUMP_OFF_1/off_on_timer_0/count[1]  (.D(
        \DUMP_OFF_1/off_on_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/count_4[1] ));
    DFN1E0 \DDS_0/dds_state_0/para[34]  (.D(
        \DDS_0/dds_state_0/para_9[34] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[34]_net_1 ));
    OR2 \top_code_0/s_acqnum_1_sqmuxa_0_o2  (.A(\top_code_0/N_142 ), 
        .B(\xa_c[4] ), .Y(\top_code_0/N_150 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m46_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[13] ));
    OR2A \top_code_0/relay_close_1_sqmuxa_0_o2_0  (.A(\xa_c[0] ), .B(
        \xa_c[1] ), .Y(\top_code_0/N_147 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[8]  (.A(
        \scalestate_0/s_acqnum_7[8] ), .B(\scalestate_0_s_acqnum[8] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_555 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i6_mux ));
    DFN1 \DUMP_ON_0/off_on_timer_0/count[2]  (.D(
        \DUMP_ON_0/off_on_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/count_5[2] ));
    DFN1E1 \noisestate_0/dectime[9]  (.D(\top_code_0_noisedata[9] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[9]_net_1 ));
    NOR3C \scalestate_0/CUTTIME180_Tini_532_e  (.A(\scalestate_0/N_66 )
        , .B(\scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 ), .C(
        \top_code_0_scalechoice_0[0] ), .Y(\scalestate_0/N_1745 ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[6]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_34_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[6] ));
    OR3 \DUMP_0/dump_coder_0/para5_RNIGBAK2[6]  (.A(
        \DUMP_0/dump_coder_0/un1_count_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_11[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_6[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[2]_net_1 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/ADD_20x20_slow_I19_Y_0 )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i4_mux ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_8  (.A(\PLUSE_0/count_2[6] ), 
        .B(\PLUSE_0/half_para[6] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[1] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m14  (.A(
        \top_code_0_n_divnum_0[5] ), .B(\top_code_0_n_divnum_0[0] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[0] ));
    AND3 \scalestate_0/necount_inc_0/AND2_1_7_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount_inc_0/inc_5_net ), .C(
        \scalestate_0/necount[6]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/Rcout_7_net ));
    DFN1 \DDS_0/dds_state_0/cs[8]  (.D(
        \DDS_0/dds_state_0/cs_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[8]_net_1 ));
    IOTRI_OR_EB \ddsfqud_pad/U0/U1  (.D(
        \DDS_0/dds_state_0/fq_ud_RNO_net_1 ), .E(VCC), .OCLK(GLA_net_1)
        , .DOUT(\ddsfqud_pad/U0/NET1 ), .EOUT(\ddsfqud_pad/U0/NET2 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_31  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[6] )
        , .B(\s_acq_change_0_s_stripnum[9] ), .C(
        \s_acq_change_0_s_stripnum[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_18  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[1] )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIE0DH[18]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[18]_net_1 ), .B(
        \sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_18[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[0]  (.A(
        \state_1ms_0_timecount[0] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_242 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m97  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_90 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_97 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[5] ));
    NOR2B \DDS_0/dds_state_0/cs_RNO[4]  (.A(
        \DDS_0/dds_state_0/cs[3]_net_1 ), .B(\DDS_0/dds_state_0/N_223 )
        , .Y(\DDS_0/dds_state_0/cs_RNO[4]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIOI4A4[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_7[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_18[0] ));
    DFN1E1 \state_1ms_0/CUTTIME[2]  (.D(\top_code_0_state_1ms_data[2] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[2]_net_1 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNO_0[11]  (.A(
        \ClockManagement_0/long_timer_0/count_c9 ), .B(
        \ClockManagement_0/long_timer_0/count[10]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c10 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIE1301[3]  (
        .A(\pd_pluse_top_0/count_6[3] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[3]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_0[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_7[0] ));
    NOR2B \ClockManagement_0/long_timer_0/clk_5K_reg2_RNO  (.A(
        \ClockManagement_0/long_timer_0/clk_5K_reg1_net_1 ), .B(net_27)
        , .Y(\ClockManagement_0/long_timer_0/clk_5K_reg2_RNO_net_1 ));
    MX2 \scalestate_0/strippluse_RNO_0[4]  (.A(
        \scalestate_0/strippluse_6[4] ), .B(
        \scalestate_0_strippluse[4] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_563 ));
    DFN1E1 \scanstate_0/dectime[10]  (.D(\top_code_0_scandata[10] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[10]_net_1 ));
    DFN1E1 \plusestate_0/PLUSETIME[11]  (.D(\top_code_0_plusedata[11] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[11]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_9  (.A(
        \timer_top_0/timer_0/N_20 ), .B(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .Y(
        \timer_top_0/timer_0/I_9_2 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[6] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[5] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_62_i ));
    NOR2A \scalestate_0/timecount_ret_88_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[10]_net_1 ), .B(\scalestate_0/N_1089 )
        , .Y(\scalestate_0/S_DUMPTIME_m[10] ));
    NOR3C \scalestate_0/ACQ180_NUM_1_sqmuxa_0_a2  (.A(
        \scalestate_0/N_67 ), .B(\top_code_0_scalechoice_0[0] ), .C(
        \scalestate_0/N_62 ), .Y(\scalestate_0/ACQ180_NUM_1_sqmuxa ));
    DFN1E1 \top_code_0/sigtimedata[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[1] ));
    MX2 \scanstate_0/timecount_1_RNO_0[6]  (.A(
        \scanstate_0/acqtime[6]_net_1 ), .B(
        \scanstate_0/dectime[6]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_64 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m28  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_29 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[4]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[30]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[31]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_516 ));
    OR3 \top_code_0/un1_state_1ms_rst_n117_47_i_o2  (.A(
        \top_code_0/N_328 ), .B(\top_code_0/N_327 ), .C(
        \top_code_0/N_330 ), .Y(\top_code_0/N_162 ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_40  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[2]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[7] ));
    DFN1 \top_code_0/scan_start_ret_2  (.D(\top_code_0/un1_xa_10 ), 
        .CLK(GLA_net_1), .Q(\top_code_0/un1_xa_10_reto ));
    DFN1 \s_acq_change_0/s_stripnum[1]  (.D(
        \s_acq_change_0/s_stripnum_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[1] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[14]_net_1 ));
    DFN1 \top_code_0/relay_close[8]  (.D(
        \top_code_0/relay_close_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[8] ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_1  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[7]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] )
        );
    MX2 \scalestate_0/strippluse_RNO_2[11]  (.A(
        \scalestate_0/STRIPNUM180_NUM[11]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[11]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_431 ));
    NOR2B \scalestate_0/CS_RNO[9]  (.A(\scalestate_0/N_1223 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO_0[9]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[0] ));
    NOR2B \DUMP_OFF_0/off_on_timer_0/count_RNO_0[4]  (.A(
        \DUMP_OFF_0/count_3[3] ), .B(
        \DUMP_OFF_0/off_on_timer_0/count_c2 ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_9_0 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/OXOR2_15_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_19_net ), 
        .B(\sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[19] ));
    NOR3C \scalestate_0/timecount_ret_35_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[9]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[9] ));
    DFN1E1 \scanstate_0/timecount_1[10]  (.D(
        \scanstate_0/timecount_5[10] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[10] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[3]  (.A(
        \s_acq_change_0/s_acqnum_5[3] ), .B(
        \s_acq_change_0_s_acqnum[3] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_73 ));
    NOR3B \DUMP_ON_0/off_on_state_0/cs_RNO[1]  (.A(OR2_2_Y), .B(
        \DUMP_ON_0/i_5[0] ), .C(\DUMP_ON_0/off_on_state_0/N_10 ), .Y(
        \DUMP_ON_0/off_on_state_0/cs_nsss[1] ));
    MX2 \scalestate_0/strippluse_RNO_2[5]  (.A(
        \scalestate_0/STRIPNUM180_NUM[5]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[5]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_425 ));
    MX2 \bri_dump_sw_0/reset_out_5  (.A(top_code_0_pluse_rst), .B(
        net_45), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/reset_out_5_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_133  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_133_Y ));
    AND2A \scalestate_0/necount_cmp_0/AND2A_0  (.A(
        \scalestate_0/necount[10]_net_1 ), .B(
        \scalestate_0/M_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/AND2A_0_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[24]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[24]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_304 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i2_mux ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m159  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_160 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[0]_net_1 ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_14  (.A(
        \scalestate_0/NE_NUM[9]_net_1 ), .B(
        \scalestate_0/necount[9]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_9 ));
    NOR2A \timer_top_0/state_switch_0/state_start5_0_0_a2_2_0  (.A(
        top_code_0_noise_start), .B(top_code_0_scan_start), .Y(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_2_0_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_63  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_63_Y ));
    NOR3C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en_net_1 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_11 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_1_sqmuxa ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]  
        (.D(\s_acq_change_0_s_acqnum[12] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]_net_1 )
        );
    DFN1 \DDS_0/dds_timer_0/count[1]  (.D(\DDS_0/dds_timer_0/count_n1 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[1] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m298  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_299 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[5]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[5] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[5] ));
    NOR2B \scalestate_0/timecount_ret_8_RNO_3  (.A(
        \scalestate_0/OPENTIME[3]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[3] ));
    NOR3C \scalestate_0/OPENTIME_TEL_576_e  (.A(\scalestate_0/N_64 ), 
        .B(\scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0_0[0] ), 
        .Y(\scalestate_0/N_1789 ));
    DFN1 \timer_top_0/timer_0/timedata[14]  (.D(
        \timer_top_0/timer_0/timedata_4[14] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[14]_net_1 ));
    DFN1E1 \noisestate_0/dectime[6]  (.D(\top_code_0_noisedata[6] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[6]_net_1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[11]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c10 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n11 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m285  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_284 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_285 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_286 ));
    MX2 \scanstate_0/timecount_1_RNO_0[11]  (.A(
        \scanstate_0/dectime[11]_net_1 ), .B(
        \scanstate_0/acqtime[11]_net_1 ), .S(\scanstate_0/CS[4]_net_1 )
        , .Y(\scanstate_0/N_69 ));
    XO1 \DUMP_0/dump_coder_0/para3_RNIM0V21[2]  (.A(
        \DUMP_0/count_1[2] ), .B(\DUMP_0/dump_coder_0/para3[2]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_2_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_3[0] ));
    OA1B \plusestate_0/CS_RNO[2]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[2]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[2] )
        , .Y(\plusestate_0/CS_RNO_0[2]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[2]  (.D(\top_code_0_scaledatain[2] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[2]_net_1 ));
    DFN1 \bri_dump_sw_0/reset_out  (.D(
        \bri_dump_sw_0/reset_out_0_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_reset_out));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i20_mux ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[10]  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n10 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i22_mux ));
    DFN1E1 \scalestate_0/DUMPTIME[9]  (.D(\top_code_0_scaledatain[9] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[9]_net_1 ));
    MX2 \scalestate_0/CS_RNO_0[17]  (.A(\scalestate_0/CS[17]_net_1 ), 
        .B(\scalestate_0/CS[16]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1230 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m44_4 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_52_i ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[5]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n5 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ));
    DFN1E1 \scalestate_0/DUMPTIME[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[14]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[5]  (.D(
        \DUMP_0/dump_coder_0/para4_4[5]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[5]_net_1 ));
    AO1A \scalestate_0/timecount_ret_7_RNI68SS  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .B(
        \scalestate_0/timecount_cnst_m_0_reto[3] ), .C(
        \scalestate_0/timecount_20_iv_10_reto[3] ), .Y(
        \scalestate_0_timecount[3] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIOTRO1[11]  (.A(
        \sd_acq_top_0/count_1[11] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[11]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_12[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_3[0] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[12]  (.D(
        \top_code_0_dds_configdata[11] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[12]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[3] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNITI8D[14]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[14]_net_1 )
        , .B(\pd_pluse_top_0/count[14] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_14[0] ));
    NOR2A \s_acq_change_0/s_acqnum_RNO_1[14]  (.A(
        \top_code_0_s_acqnum_2[14] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[14] ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[10]  (.D(
        \DUMP_0/dump_coder_0/para4_4[10]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[10]_net_1 ));
    DFN1 \DDS_0/dds_state_0/cs[6]  (.D(
        \DDS_0/dds_state_0/cs_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[6]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_choice[2]  (.D(\GPMI_0_dataout[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_choice_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_choice[2] ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNII3T21[13]  
        (.A(\pd_pluse_top_0/count[13] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[13]_net_1 ), 
        .C(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_10[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_2[0] ));
    NOR2B \ClockManagement_0/clk_div500_0/un1_count_1_I_44  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_TMP[0] ), .B(
        \ClockManagement_0/clk_div500_0/count[1]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_1[0] ));
    DFN1E1 \scanstate_0/timecount_1[5]  (.D(
        \scanstate_0/timecount_5[5] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[5] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[11]  (.A(
        \scalestate_0/ACQ180_NUM[11]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[11]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_459 ));
    DFN1 \state_1ms_0/timecount[3]  (.D(
        \state_1ms_0/timecount_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[3] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIUN1G[5]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[5]_net_1 ), 
        .B(\pd_pluse_top_0/count_1[5] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_5[0] ));
    OA1B \noisestate_0/CS_RNO[3]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[3]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[3] )
        , .Y(\noisestate_0/CS_RNO[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_1_Y ));
    OA1B \plusestate_0/CS_RNO[6]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[6]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[6] )
        , .Y(\plusestate_0/CS_RNO_0[6]_net_1 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[20]  (.A(
        \DDS_0/dds_state_0/N_468 ), .B(\DDS_0/dds_state_0/N_467 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[20] ), .Y(
        \DDS_0/dds_state_0/N_123 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[5]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[5] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_3[5] ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNIHKCG[5]  (.A(
        \DUMP_0/dump_coder_0/para2[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_5[0] ));
    DFN1 \DUMP_OFF_1/off_on_state_0/cs[0]  (.D(
        \DUMP_OFF_1/off_on_state_0/N_36_i ), .CLK(GLA_net_1), .Q(
        DUMP_OFF_1_dump_off));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m216  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[9] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_217 ));
    DFN1 \scalestate_0/CS[8]  (.D(\scalestate_0/CS_RNO_0[8]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[8]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m291  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_292 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[5] ));
    MX2B \plusestate_0/timecount_1_RNO[5]  (.A(\plusestate_0/N_76 ), 
        .B(\plusestate_0/N_251 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[5] ));
    NOR2B \scalestate_0/timecount_ret_68_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[14]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[14] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[32]  (.D(
        \top_code_0_dds_configdata[15] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[32]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO[12]  (.A(\state_1ms_0/N_79 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_10  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_10_Y ));
    MX2 \scalestate_0/necount_RNO_0[5]  (.A(\scalestate_0/necount1[5] )
        , .B(\scalestate_0/necount[5]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_735 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_77  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_163_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_157_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_77_Y ));
    DFN1P0 \PLUSE_0/bri_state_0/cs[0]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[0] ), .CLK(ddsclkout_c), .PRE(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[0]_net_1 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[1]  (.D(\top_code_0_scaledatain[1] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[1]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/state_start5_0_0_a2_0  (.A(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_0_0 ), .B(
        \timer_top_0/state_switch_0/N_284 ), .Y(
        \timer_top_0/state_switch_0/N_168 ));
    DFN1E1 \plusestate_0/timecount_1[6]  (.D(
        \plusestate_0/timecount_5[6] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[6] ));
    NOR2B \top_code_0/state_1ms_start_ret_1_RNIRKNJ1  (.A(
        \top_code_0/N_795_reto ), .B(\top_code_0/net_27_reto ), .Y(
        top_code_0_state_1ms_start));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_50_i ));
    NOR2B 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNI9ND34[9]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c8 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c9 ));
    NOR2B \top_code_0/un1_xa_10_0_a2_2  (.A(\top_code_0/N_337 ), .B(
        \top_code_0/N_336 ), .Y(\top_code_0/un1_xa_10_2 ));
    OA1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_86  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_23_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_126_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_86_Y ));
    MX2B \scanstate_0/timecount_1_RNO[0]  (.A(\scanstate_0/N_58 ), .B(
        net_33_0), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[0] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_2  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m38 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[4] )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_35  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_26_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_109_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_35_Y ));
    NOR3C \scalestate_0/CUTTIME90_488_e  (.A(\scalestate_0/N_62 ), .B(
        \scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/N_1701 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_39  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_53_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_8_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_39_Y ));
    NOR3C \state_1ms_0/S_DUMPTIME_1_sqmuxa_0_a2  (.A(
        \top_code_0_state_1ms_lc[0] ), .B(\top_code_0_state_1ms_lc[1] )
        , .C(\state_1ms_0/N_17 ), .Y(\state_1ms_0/S_DUMPTIME_1_sqmuxa )
        );
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_50_i ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[20]  (.D(
        \top_code_0_dds_configdata[3] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[20]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[4]  (.D(
        \DUMP_0/dump_coder_0/para2_4[4]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[4]_net_1 ));
    OR3 \scalestate_0/timecount_ret_8_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[3] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[3] ), .C(
        \scalestate_0/timecount_20_iv_2[3] ), .Y(
        \scalestate_0/timecount_20_iv_7[3] ));
    MX2 \state_1ms_0/timecount_RNO_0[9]  (.A(
        \state_1ms_0/timecount_8[9] ), .B(\state_1ms_0_timecount[9] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_76 ));
    NOR3B \DUMP_0/dump_state_0/cs_RNO_0[5]  (.A(
        \DUMP_0/dump_state_0/N_206 ), .B(\DUMP_0/dump_state_0/N_167 ), 
        .C(\DUMP_0/dump_state_0/cs[4]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_193 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_72  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_72_Y ));
    DFN1E1 \plusestate_0/timecount_1[1]  (.D(
        \plusestate_0/timecount_5[1] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[1] ));
    OR3 \scalestate_0/timecount_ret_RNO  (.A(\scalestate_0/N_1197 ), 
        .B(\scalestate_0/CS[16]_net_1 ), .C(\scalestate_0/N_1206 ), .Y(
        \scalestate_0/timecount_cnst[5] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m43_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] ));
    NOR2A \scalestate_0/timecount_ret_53_RNO_3  (.A(
        \scalestate_0/CUTTIME90[18]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[18] ));
    DFN1 \plusestate_0/soft_d  (.D(\plusestate_0/soft_d_RNO_1_net_1 ), 
        .CLK(GLA_net_1), .Q(plusestate_0_soft_d));
    NOR2B \scalestate_0/CS_RNO[5]  (.A(\scalestate_0/N_1220 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO_1[5] ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[8]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[8]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/i_0[8] ));
    IOTRI_OB_EB \syn_md_out_pad/U0/U1  (.D(syn_md_out_c), .E(VCC), 
        .DOUT(\syn_md_out_pad/U0/NET1 ), .EOUT(
        \syn_md_out_pad/U0/NET2 ));
    OA1A \PLUSE_0/bri_coder_0/half_0_I_23  (.A(
        \PLUSE_0/bri_coder_0/N_6 ), .B(\PLUSE_0/bri_coder_0/N_8 ), .C(
        \PLUSE_0/bri_coder_0/N_7 ), .Y(\PLUSE_0/bri_coder_0/N_11 ));
    NOR2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y ));
    NOR2B \DUMP_0/dump_timer_0/count_RNI25BE1[3]  (.A(
        \DUMP_0/dump_timer_0/count_c2 ), .B(\DUMP_0/count_1[3] ), .Y(
        \DUMP_0/dump_timer_0/count_c3 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[11] ));
    MX2 \nsctrl_choice_0/intertodsp_RNO_0  (.A(
        scanstate_0_state_over_n), .B(noisestate_0_state_over_n), .S(
        top_code_0_n_s_ctrl_0), .Y(\nsctrl_choice_0/intertodsp_5 ));
    DFN1 \state_1ms_0/timecount[11]  (.D(
        \state_1ms_0/timecount_RNO[11]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[11] ));
    NOR2B \DUMP_OFF_1/off_on_timer_0/count_RNO_0[4]  (.A(
        \DUMP_OFF_1/count_4[3] ), .B(
        \DUMP_OFF_1/off_on_timer_0/count_c2 ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_9_0 ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_10  (.A(
        \timer_top_0/dataout[5] ), .B(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_10_Y ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i12_mux ));
    DFN1 \DUMP_0/dump_coder_0/i[1]  (.D(
        \DUMP_0/dump_coder_0/i_RNO_0[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_2[1] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[7]  (.D(
        \top_code_0_state_1ms_data[7] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[7]_net_1 ));
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_36  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[0] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[1] ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[2] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[3] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m118  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_117 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_118 ), .S(
        \top_code_0_s_addchoice_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_119 ));
    IOIN_IB \xa_pad[18]/U0/U1  (.YIN(\xa_pad[18]/U0/NET1 ), .Y(
        \xa_c[18] ));
    NOR2B \top_code_0/dump_sustain_RNO  (.A(\top_code_0/N_808 ), .B(
        net_27), .Y(\top_code_0/dump_sustain_RNO_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[14]_net_1 ));
    AND3 \PLUSE_0/bri_coder_0/half_0_I_4  (.A(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[2] ), .B(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[1] ), .C(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[0] ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[1] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[10]  (.A(
        \timer_top_0/state_switch_0/N_252 ), .B(
        \timer_top_0/state_switch_0/N_254 ), .C(
        \timer_top_0/state_switch_0/N_253 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[10] ));
    MX2C \DUMP_OFF_1/off_on_state_0/cs_RNO_0[1]  (.A(
        \DUMP_OFF_1/off_on_state_0/cs[1]_net_1 ), .B(
        \DUMP_OFF_1/i_4[1] ), .S(DUMP_OFF_1_dump_off), .Y(
        \DUMP_OFF_1/off_on_state_0/N_10 ));
    DFN1E1 \top_code_0/s_addchoice_5[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_5[4] ));
    DFN1 \state_1ms_0/timecount[18]  (.D(
        \state_1ms_0/timecount_RNO[18]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[18] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_41_i ));
    MX2B \scanstate_0/timecount_1_RNO[11]  (.A(\scanstate_0/N_69 ), .B(
        \scanstate_0/N_196 ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[11] ));
    DFN1 \state_1ms_0/timecount[12]  (.D(
        \state_1ms_0/timecount_RNO[12]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[12] ));
    OR3A \scalestate_0/timecount_ret_17_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/N_258_0 ), .C(
        \scalestate_0/un1_timecount_2_sqmuxa_4 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[0]  (.D(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_6[0] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/i_6[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_146  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_146_Y ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n2 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        );
    XOR2 \PLUSE_0/bri_timer_0/count_RNO[0]  (.A(\PLUSE_0/count_8[0] ), 
        .B(\PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count_e0 ));
    AO1 \DDS_0/dds_state_0/para_RNO[33]  (.A(
        \DDS_0/dds_state_0/para[33]_net_1 ), .B(
        \DDS_0/dds_state_0/N_538_0 ), .C(\DDS_0/dds_state_0/N_522 ), 
        .Y(\DDS_0/dds_state_0/para_9[33] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i14_mux ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[4]  (.D(
        \DUMP_0/dump_coder_0/para4_4[4]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[4]_net_1 ));
    AOI1B \DDS_0/dds_state_0/cs_RNO[2]  (.A(\DDS_0/dds_state_0/N_228 ), 
        .B(\DDS_0/dds_state_0/N_225 ), .C(\DDS_0/dds_state_0/N_223 ), 
        .Y(\DDS_0/dds_state_0/N_38 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[12]  (.D(
        \top_code_0_state_1ms_data[12] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[12]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m94  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_95 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i2_mux ));
    OR3 \scalestate_0/fst_lst_pulse_RNO_1  (.A(
        \scalestate_0/fst_lst_pulse8_NE_4 ), .B(
        \scalestate_0/fst_lst_pulse8_NE_3 ), .C(
        \scalestate_0/fst_lst_pulse8_NE_8 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[14]  (.A(
        \plusestate_0_timecount[14] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_264 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[7]_net_1 ));
    DFN1 \state_1ms_0/CS_i[0]  (.D(\state_1ms_0/CS_i_RNO_1[0] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS_i[0]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[14]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[14] ), .CLK(ddsclkout_c)
        , .Q(\sd_acq_top_0/sd_sacq_state_0/cs[14]_net_1 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[2]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[2] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[2]_net_1 ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_1_5_inst  (.A(
        \scalestate_0/necount_inc_0/Rcout_7_net ), .B(
        \scalestate_0/necount[7]_net_1 ), .Y(
        \scalestate_0/necount1[7] ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNICA8P[10]  (.A(
        \DUMP_0/dump_coder_0/para5[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_10[0] ));
    IOTRI_OB_EB \relay_close_pad[9]/U0/U1  (.D(\relay_close_c[9] ), .E(
        VCC), .DOUT(\relay_close_pad[9]/U0/NET1 ), .EOUT(
        \relay_close_pad[9]/U0/NET2 ));
    OA1B \noisestate_0/CS_RNO[5]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[5]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[5] )
        , .Y(\noisestate_0/CS_RNO[5]_net_1 ));
    MX2 \top_code_0/noise_start_ret_2_RNI09J61  (.A(
        \top_code_0/top_code_0_noise_start_reto ), .B(
        \top_code_0/un1_xa_13_reto ), .S(\top_code_0/N_114_reto ), .Y(
        \top_code_0/N_799_reto ));
    OR3 \state_1ms_0/timecount_RNO_1[2]  (.A(
        \state_1ms_0/timecount_8_iv_1[2] ), .B(
        \state_1ms_0/timecount_8_iv_0[2] ), .C(
        \state_1ms_0/timecount_8_iv_2[2] ), .Y(
        \state_1ms_0/timecount_8_iv[2] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[0] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/dataout[13]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[13] ), .B(
        top_code_0_n_s_ctrl_1), .Y(\Signal_Noise_Acq_0_dataout[13] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m7  
        (.A(\s_acq_change_0_s_stripnum[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[2]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i4_mux ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIT5QK[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_11[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[19]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[19]_net_1 ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_5  (.A(
        \scalestate_0/NE_NUM[10]_net_1 ), .B(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_10 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[5]  (.A(
        \top_code_0_s_acqnum_2[5] ), .B(\scalestate_0_s_acqnum[5] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[5] ));
    XA1A \CAL_0/cal_div_0/cal_RNO_0  (.A(\CAL_0/cal_div_0/clear_n ), 
        .B(cal_out_c), .C(scanstate_0_calctrl), .Y(
        \CAL_0/cal_div_0/N_35 ));
    NOR2A \top_code_0/cal_data_1_sqmuxa_0_a2_1  (.A(net_27), .B(
        \top_code_0/N_165 ), .Y(\top_code_0/cal_data_1_sqmuxa_1 ));
    NOR2A \DUMP_OFF_0/off_on_timer_0/count_RNO[0]  (.A(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_OFF_0/count_3[0] ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_n0 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_8  (.A(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[2]_net_1 ), .Y(
        \timer_top_0/timer_0/N_20 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_3  (.A(\ADC_c[7] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ));
    OR3 \DUMP_0/dump_coder_0/para2_RNI44SD2[6]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_3_11[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_3_NE_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_6[0] ));
    MX2 \scalestate_0/strippluse_RNO_0[9]  (.A(
        \scalestate_0/strippluse_6[9] ), .B(
        \scalestate_0_strippluse[9] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_568 ));
    DFN1E0 \DDS_0/dds_state_0/para[15]  (.D(\DDS_0/dds_state_0/N_159 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[15]_net_1 ));
    OR3A \top_code_0/acqclken_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_164 ), .Y(
        \top_code_0/N_199 ));
    DFN1 \scalestate_0/s_acq180  (.D(\scalestate_0/s_acq180_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(s_acq180_c));
    IOTRI_OB_EB \Q3Q6_pad/U0/U1  (.D(Q3Q6_c), .E(VCC), .DOUT(
        \Q3Q6_pad/U0/NET1 ), .EOUT(\Q3Q6_pad/U0/NET2 ));
    MX2A \state_1ms_0/timecount_RNO_0[2]  (.A(
        \state_1ms_0/timecount_8_iv[2] ), .B(
        \state_1ms_0_timecount[2] ), .S(\state_1ms_0/CS[9]_net_1 ), .Y(
        \state_1ms_0/N_69 ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_5  (.A(
        \scalestate_0/necount[7]_net_1 ), .B(
        \scalestate_0/NE_NUM[7]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_5_Y ));
    DFN1E1 \top_code_0/pd_pluse_data[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[15] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_0  (.A(
        \scalestate_0/NE_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_0_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_88  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_88_Y ));
    OR2 \PLUSE_0/qq_coder_0/i_reg10_NE[0]  (.A(
        \PLUSE_0/qq_coder_0/i_reg10_NE_3[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_0/i_reg10_NE_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_NE[0]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[15]_net_1 ));
    DFN1 \plusestate_0/CS[2]  (.D(\plusestate_0/CS_RNO_0[2]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[2]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_138  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_19_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_99_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_138_Y ));
    DFN1 \scalestate_0/strippluse[4]  (.D(
        \scalestate_0/strippluse_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[4] ));
    IOIN_IB \zcs2_pad/U0/U1  (.YIN(\zcs2_pad/U0/NET1 ), .Y(zcs2_c));
    OR3 \scalestate_0/timecount_ret_68_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[14] ), .B(
        \scalestate_0/OPENTIME_TEL_m[14] ), .C(
        \scalestate_0/timecount_20_iv_4[14] ), .Y(
        \scalestate_0/timecount_20_iv_8[14] ));
    DFN1E0 \DDS_0/dds_state_0/para[11]  (.D(\DDS_0/dds_state_0/N_87 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[11]_net_1 ));
    IOIN_IB \xa_pad[8]/U0/U1  (.YIN(\xa_pad[8]/U0/NET1 ), .Y(\xa_c[8] )
        );
    OR3 \topctrlchange_0/interupt_RNO_1  (.A(
        \topctrlchange_0/interin2_m ), .B(\topctrlchange_0/interin3_m )
        , .C(\topctrlchange_0/interin1_m ), .Y(
        \topctrlchange_0/un1_interin1[0] ));
    NOR3C \DUMP_OFF_1/off_on_state_0/cs_RNO[0]  (.A(
        nsctrl_choice_0_dumponoff_rst), .B(\DUMP_OFF_1/i_4[0] ), .C(
        \DUMP_OFF_1/off_on_state_0/N_42_i ), .Y(
        \DUMP_OFF_1/off_on_state_0/N_36_i ));
    XA1 \DDS_0/dds_timer_0/count_RNO[5]  (.A(
        \DDS_0/dds_timer_0/count_c4 ), .B(\DDS_0/count[5] ), .C(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DDS_0/dds_timer_0/count_n5 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[10]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[10] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_0[10] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_0_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_0_net ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[9]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[9] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_1[9] ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg_RNIS2Q11[3]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[3]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_2 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[1]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_i ), 
        .C(\s_acq_change_0_s_stripnum[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i2_mux ));
    AO1C \noisestate_0/CS_RNO_0[6]  (.A(\noisestate_0/CS[5]_net_1 ), 
        .B(timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[6] ));
    NOR2B \DUMP_0/dump_timer_0/count_RNI8AO21[2]  (.A(
        \DUMP_0/dump_timer_0/count_c1 ), .B(\DUMP_0/count_1[2] ), .Y(
        \DUMP_0/dump_timer_0/count_c2 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_5_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_5_net ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[9]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[9]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/i[9] ));
    NOR2B \scalestate_0/timecount_ret_55_RNO  (.A(
        \scalestate_0/OPENTIME_TEL[19]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[19] ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[7]_net_1 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[8]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[8] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[8]_net_1 ));
    DFN1 \scalestate_0/CS[21]  (.D(\scalestate_0/CS_RNO[21]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[21]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m301  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_298 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_301 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_302 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_10_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_44_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_81_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_10_inst ));
    NOR2A \scalestate_0/timecount_ret_82_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[4]_net_1 ), .B(\scalestate_0/N_1089 ), 
        .Y(\scalestate_0/S_DUMPTIME_m[4] ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[8]  (.D(
        \DUMP_0/dump_coder_0/para4_4[8]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[8]_net_1 ));
    MX2 \plusestate_0/timecount_1_RNO_0[3]  (.A(
        \plusestate_0/DUMPTIME[3]_net_1 ), .B(
        \plusestate_0/PLUSETIME[3]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_74 ));
    MX2 \PLUSE_0/bri_timer_0/count[3]/U0  (.A(\PLUSE_0/count_8[3] ), 
        .B(\PLUSE_0/bri_timer_0/count_n3 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[3]/Y ));
    OR3 \PLUSE_0/bri_state_0/up_RNO  (.A(\PLUSE_0/bri_state_0/N_144 ), 
        .B(\PLUSE_0/bri_state_0/cs[3]_net_1 ), .C(
        \PLUSE_0/bri_state_0/N_178 ), .Y(\PLUSE_0/bri_state_0/down30 ));
    AND3B \top_code_0/un1_state_1ms_rst_n117_3_i_a2  (.A(
        \top_code_0/N_161 ), .B(\top_code_0/N_171 ), .C(
        \top_code_0/N_332 ), .Y(\top_code_0/N_259 ));
    DFN1E1 \top_code_0/bri_datain[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[2] ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/FOR2_8_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_10_net ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[10] ));
    NOR2A \scalestate_0/timecount_ret_64_RNO_0  (.A(
        \scalestate_0/ACQTIME[13]_net_1 ), .B(\scalestate_0/N_1065 ), 
        .Y(\scalestate_0/ACQTIME_m[13] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[18]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[19]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_504 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[9]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_26_0 ), .Y(
        \timer_top_0/timer_0/timedata_4[9] ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[10]  (.A(
        \top_code_0_dumpdata_0[10] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[10]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_6[3]  (.A(
        \DUMP_0/dump_coder_0/para1[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_3[0] ));
    OA1B \state_1ms_0/CS_RNO[5]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[5]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[5] ), 
        .Y(\state_1ms_0/CS_RNO_3[5] ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BFF1_3_inst  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_3_net ));
    DFN1 \plusestate_0/sw_acq1  (.D(\plusestate_0/sw_acq1_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(plusestate_0_sw_acq1));
    DFN1E1 \top_code_0/n_load  (.D(\top_code_0/N_72 ), .CLK(GLA_net_1), 
        .E(net_27), .Q(top_code_0_n_load));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_2_i ));
    DFN1E1 \scalestate_0/timecount_ret_28  (.D(
        \scalestate_0/timecount_20_iv_9[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_9_reto[1] ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_1_5_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_7_net ), 
        .B(\sd_acq_top_0/count_3[7] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[7] ));
    OR2B \scanstate_0/CS_RNICADM[4]  (.A(\scanstate_0/CS[4]_net_1 ), 
        .B(net_33), .Y(\scanstate_0/N_194 ));
    XA1 \DUMP_OFF_0/off_on_timer_0/count_RNO[4]  (.A(
        \DUMP_OFF_0/off_on_timer_0/count_9_0 ), .B(
        \DUMP_OFF_0/count_3[4] ), .C(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_n4 ));
    DFN0 \DSTimer_0/DFN0_0  (.D(top_code_0_dump_sustain), .CLK(
        GLA_net_1), .Q(\DSTimer_0/net_0 ));
    DFN1E1 \scanstate_0/timecount_1[7]  (.D(
        \scanstate_0/timecount_5[7] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[7] ));
    NOR3C \scalestate_0/CUTTIMEI90_554_e  (.A(\scalestate_0/N_64 ), .B(
        \scalestate_0/N_65 ), .C(\top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/N_1767 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/en  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/en_RNO_net_1 ), .CLK(
        ddsclkout_c), .Q(pd_pulse_en_c));
    AO1 \scalestate_0/timecount_ret_69_RNO_2  (.A(
        \scalestate_0/CUTTIME180_TEL[15]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[15] )
        , .Y(\scalestate_0/timecount_20_iv_3[15] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[5]  (.D(
        \top_code_0_pd_pluse_data[5] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[5]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[10]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[11]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_293 ));
    OR2A \top_code_0/scale_rst_0_0_RNI25ID3  (.A(net_27), .B(
        \top_code_0/N_801 ), .Y(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ));
    DFN1E1 \scalestate_0/PLUSETIME90[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[14]_net_1 ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[10]  (.A(
        \PLUSE_0/bri_state_0/cs[10]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs[9]_net_1 ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_0[10] ));
    AO1C \DUMP_0/dump_coder_0/un1_para114_6  (.A(
        \DUMP_0/dump_coder_0/para15_net_1 ), .B(
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ), .C(
        top_code_0_dumpload), .Y(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/YAND2B_22_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_5_net ), 
        .C(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[17]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[17]_net_1 ));
    OR3 \top_code_0/nstateload_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_149 ), .Y(
        \top_code_0/N_211 ));
    MX2 \scalestate_0/CS_RNO_0[14]  (.A(\scalestate_0/CS[14]_net_1 ), 
        .B(\scalestate_0/CS[13]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1227 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[31]  (.A(
        \DDS_0/dds_state_0/N_569 ), .B(\top_code_0_dds_configdata[14] )
        , .Y(\DDS_0/dds_state_0/N_517 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIUQJO3[14]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_3[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_2[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_17[0] ));
    AO1B \scalestate_0/CS_RNIDSG82[18]  (.A(\scalestate_0/N_1310 ), .B(
        timer_top_0_clk_en_scale), .C(top_code_0_scale_rst_1), .Y(
        \scalestate_0/un1_CS6_33 ));
    DFN1 \timer_top_0/state_switch_0/dataout[0]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[0]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m86  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_87 ));
    OR3 \DUMP_0/dump_coder_0/para4_RNICUQC2[11]  (.A(
        \DUMP_0/dump_coder_0/un1_count_1_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_11[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_1_NE_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_6[0] ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_5  (.A(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .B(
        \timer_top_0/dataout[20] ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_9_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_5_Y ));
    NOR2B \state_1ms_0/timecount_RNO_3[10]  (.A(
        \state_1ms_0/CUTTIME[10]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[10] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[0]_net_1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[7]  (.A(
        \s_acq_change_0/s_stripnum_5[7] ), .B(
        \s_acq_change_0_s_stripnum[7] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_63 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i2_mux ));
    NOR3 \DDS_0/dds_state_0/para_RNO[32]  (.A(
        \DDS_0/dds_state_0/N_314 ), .B(\DDS_0/dds_state_0/N_313 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[32] ), .Y(
        \DDS_0/dds_state_0/N_27 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[6]  (.A(
        \timer_top_0/state_switch_0/N_210 ), .B(
        \timer_top_0/state_switch_0/N_211 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[6] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[6]_net_1 ));
    RAM512X18 #( .MEMORYFILE("RAM_R1C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R1C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_1_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_1_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_0_net ));
    AND3 \CAL_0/cal_div_0/un3_count_I_10  (.A(
        \CAL_0/cal_div_0/count[0]_net_1 ), .B(
        \CAL_0/cal_div_0/count[1]_net_1 ), .C(
        \CAL_0/cal_div_0/count[2]_net_1 ), .Y(
        \CAL_0/cal_div_0/DWACT_FINC_E[0] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[6]  (.A(\scalestate_0/N_454 ), 
        .B(\scalestate_0/ACQECHO_NUM[6]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[6] ));
    DFN1E0 \DDS_0/dds_state_0/para[6]  (.D(\DDS_0/dds_state_0/N_44 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[6]_net_1 ));
    IOPAD_BI \xd_pad[4]/U0/U0  (.D(\xd_pad[4]/U0/NET1 ), .E(
        \xd_pad[4]/U0/NET2 ), .Y(\xd_pad[4]/U0/NET3 ), .PAD(xd[4]));
    AO1 \scalestate_0/timecount_ret_65_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[13]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[13] ), .Y(
        \scalestate_0/timecount_20_iv_4[13] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_6_inst  (.A(
        \sd_acq_top_0/count_10[3] ), .B(\sd_acq_top_0/count_10[4] ), 
        .C(\sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ));
    OR3 \scalestate_0/M_pulse_RNO_4  (.A(\scalestate_0/M_pulse8_NE_2 ), 
        .B(\scalestate_0/M_pulse8_NE_1 ), .C(
        \scalestate_0/M_pulse8_NE_5 ), .Y(\scalestate_0/M_pulse8_NE_8 )
        );
    DFN1E1 \noisestate_0/acqtime[0]  (.D(\top_code_0_noisedata[0] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[0]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[19]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[19]_net_1 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_56  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_56_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_5_0 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[1]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n1 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0  
        (.A(\top_code_0_sd_sacq_choice[2] ), .B(
        top_code_0_sd_sacq_load), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 )
        );
    DFN1E1 \scanstate_0/acqtime[11]  (.D(\top_code_0_scandata[11] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[11]_net_1 ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIE9EO1[7]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_10[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_13[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_3[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_9[0] ));
    DFN1E1 \scalestate_0/S_DUMPTIME[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[6]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[11]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i14_mux ));
    OR3 \top_code_0/state_1ms_load_RNO_0  (.A(\top_code_0/N_152 ), .B(
        \top_code_0/N_163 ), .C(\top_code_0/N_159 ), .Y(
        \top_code_0/N_197 ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[0]  (.A(\scalestate_0/N_547 ), 
        .B(top_code_0_scale_rst_5), .Y(
        \scalestate_0/s_acqnum_1_RNO[0]_net_1 ));
    OR3 \PLUSE_0/qq_coder_1/i_reg10_NE_3[0]  (.A(
        \PLUSE_0/qq_coder_1/i_reg10_2[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_1/i_reg10_3[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_1/i_reg10_NE_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_NE_3[0]_net_1 ));
    DFN1 \scalestate_0/s_acqnum_1[7]  (.D(
        \scalestate_0/s_acqnum_1_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[7] ));
    DFN1E1 \top_code_0/scaledatain[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[11] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_3_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_68_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_35_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_3_inst ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[14]_net_1 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ));
    DFN1E1 \scalestate_0/M_NUM[8]  (.D(\top_code_0_scaledatain[8] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[8]_net_1 ));
    AO1A \timer_top_0/state_switch_0/state_over_n_RNO_2  (.A(
        plusestate_0_state_over_n), .B(
        \timer_top_0/state_switch_0/N_297 ), .C(
        \timer_top_0/state_switch_0/N_280 ), .Y(
        \timer_top_0/state_switch_0/state_over_n_0_i_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_64_i ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_19  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] )
        , .C(\s_acq_change_0_s_stripnum[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7 ));
    NOR2B \top_code_0/relay_on_RNO[9]  (.A(\top_code_0/N_818 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[9]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[18]  (.D(\top_code_0_scaledatain[2] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1681 ), .Q(
        \scalestate_0/OPENTIME[18]_net_1 ));
    XA1C \DSTimer_0/dump_sustain_timer_0/start_RNO_1  (.A(
        \DSTimer_0/dump_sustain_timer_0/count[2]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/data[2]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/un1_data_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/start11_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i12_mux ));
    DFN1E1 \top_code_0/s_addchoice_0[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_0[2] ));
    DFN1E1 \scanstate_0/dectime[7]  (.D(\top_code_0_scandata[7] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[7]_net_1 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[6]  (.A(
        \scalestate_0/s_acqnum_7[6] ), .B(\scalestate_0_s_acqnum[6] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_553 ));
    AO1 \state_1ms_0/timecount_RNO_2[9]  (.A(
        \state_1ms_0/M_DUMPTIME[9]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[9] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[9] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i12_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[19]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[19]_net_1 ));
    MX2 \scalestate_0/strippluse_RNO_2[2]  (.A(
        \scalestate_0/STRIPNUM180_NUM[2]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[2]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_422 ));
    DFN1C0 \PLUSE_0/bri_coder_0/i[4]/U1  (.D(
        \PLUSE_0/bri_coder_0/i[4]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/i_1[4] ));
    NOR3C \CAL_0/cal_div_0/count_RNO[5]  (.A(net_33_0), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(\CAL_0/cal_div_0/I_14 ), 
        .Y(\CAL_0/cal_div_0/count_5[5] ));
    NOR3C \scalestate_0/timecount_ret_47_RNO_1  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[16]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[16] ));
    DFN1E0 \DDS_0/dds_state_0/para[29]  (.D(\DDS_0/dds_state_0/N_131 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[29]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_3[7]  (.A(
        \state_1ms_0/CUTTIME[7]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[7] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[0]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[4]_net_1 ));
    MX2 \scalestate_0/CS_RNO_0[19]  (.A(\scalestate_0/CS[19]_net_1 ), 
        .B(\scalestate_0/CS[3]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1231 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_9  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_9_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[14]_net_1 ));
    DFN1E1 \top_code_0/bri_datain[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[6] ));
    MX2 \top_code_0/relay_on_RNO_0[4]  (.A(\relay_on_c[4] ), .B(
        \GPMI_0_dataout[4] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_813 ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_2_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(\pd_pluse_top_0/count_6[3] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[3] ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIAFFH[1]  (.A(
        \DUMP_0/dump_coder_0/para3[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_1[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_141  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_141_Y ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[2]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[2] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[11] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[4]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n4 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[16]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[17]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_297 ));
    NOR2B \scalestate_0/necount_RNO[3]  (.A(\scalestate_0/N_733 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[3]_net_1 ));
    AND3B \pd_pluse_top_0/pd_pluse_state_0/cs_RNIO7AQ[11]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[11]_net_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[12]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_srsts_0_i_a5_1[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_195 ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIDOOK[1]  (.A(
        \DUMP_0/dump_coder_0/para6[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_1[0] ));
    DFN1E0 \DDS_0/dds_state_0/para[10]  (.D(\DDS_0/dds_state_0/N_16 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[10]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m52  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[0] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_53 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[9]  (.D(
        \top_code_0_pd_pluse_data[9] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[9]_net_1 ));
    XA1A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_13[4]  (.A(
        \pd_pluse_top_0/count[15] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[15]_net_1 ), 
        .C(net_27), .Y(\pd_pluse_top_0/pd_pluse_coder_0/i_0_0[4] ));
    AOI1 \DUMP_0/dump_state_0/cs_RNO_0[2]  (.A(
        \DUMP_0/dump_state_0/cs[1]_net_1 ), .B(\DUMP_0/i_2[1] ), .C(
        \DUMP_0/dump_state_0/cs[2]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_182 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m37  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_38_i ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[7]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[7] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[7] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[4] ));
    OA1C \scalestate_0/CS_RNIIOVH1[18]  (.A(\scalestate_0/N_1194 ), .B(
        \scalestate_0/un1_CS6_31_i_o2_0 ), .C(
        \scalestate_0/CS[18]_net_1 ), .Y(\scalestate_0/N_1310 ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[11]  (.D(
        \DUMP_0/dump_coder_0/para4_4[11]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[11]_net_1 ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_9  (.A(
        \scalestate_0/M_NUM[4]_net_1 ), .B(
        \scalestate_0/necount[4]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_9_Y ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i6_mux ));
    NOR3A \PLUSE_0/qq_state_1/cs_RNO[2]  (.A(\PLUSE_0/qq_state_1/cs4 ), 
        .B(\PLUSE_0/qq_state_1/N_89 ), .C(\PLUSE_0/qq_state_1/N_88 ), 
        .Y(\PLUSE_0/qq_state_1/cs_RNO_2[2] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m192  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_191 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_192 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_193 ));
    MX2 \scalestate_0/strippluse_RNO_0[10]  (.A(
        \scalestate_0/strippluse_6[10] ), .B(
        \scalestate_0_strippluse[10] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_569 ));
    OA1C \scalestate_0/necount_cmp_0/OA1C_0  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/M_NUM[9]_net_1 ), .C(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OA1C_0_Y ));
    DFN1 \DUMP_0/off_on_timer_1/count[3]  (.D(
        \DUMP_0/off_on_timer_1/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[3] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[20]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[20]_net_1 )
        );
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[1]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[1] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_10[1] ));
    AO1C \scalestate_0/load_out_RNO_1  (.A(\scalestate_0/un1_CS_20 ), 
        .B(\scalestate_0/un1_CS6_25_i_a3_0 ), .C(\scalestate_0/N_1196 )
        , .Y(\scalestate_0/N_1165 ));
    DFN1E1 \scalestate_0/CUTTIME180[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[7]_net_1 ));
    NOR3C \CAL_0/cal_div_0/count_RNO[4]  (.A(net_33_0), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(\CAL_0/cal_div_0/I_12 ), 
        .Y(\CAL_0/cal_div_0/count_5[4] ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_5  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_8_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_8_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_2_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_5_Y ));
    MX2 \state1ms_choice_0/soft_dump_RNO  (.A(soft_dump_net_0), .B(
        state_1ms_0_soft_dump), .S(top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/soft_dump_4 ));
    OR2A \nsctrl_choice_0/sw_acq2_RNO  (.A(net_27), .B(
        \nsctrl_choice_0/sw_acq2_5 ), .Y(
        \nsctrl_choice_0/sw_acq2_RNO_0_net_1 ));
    DFN1E1 \top_code_0/sigtimedata[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[8] ));
    OR2 \scalestate_0/timecount_ret_77_RNIE78E  (.A(
        \scalestate_0/timecount_20_iv_9_reto[6] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[6] ), .Y(
        \scalestate_0/timecount_20_iv_10_reto[6] ));
    OA1C \top_code_0/scanload_RNO  (.A(\top_code_0/N_202 ), .B(
        top_code_0_scanload), .C(\top_code_0/N_308 ), .Y(
        \top_code_0/N_100 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIUHKV[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_9[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_1[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_7[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_11[0] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m117  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[3] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_118 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i18_mux ));
    DFN1E1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[3]  
        (.D(\top_code_0_s_periodnum[3] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[3]_net_1 )
        );
    NOR3A \scalestate_0/necount_cmp_0/NOR3A_0  (.A(
        \scalestate_0/necount_cmp_0/OR2A_0_Y ), .B(
        \scalestate_0/necount_cmp_0/AO1C_2_Y ), .C(
        \scalestate_0/M_NUM[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/NOR3A_0_Y ));
    DFN1 \DUMP_OFF_1/off_on_timer_0/count[3]  (.D(
        \DUMP_OFF_1/off_on_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/count_4[3] ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_2_i ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1  (.A(\ADC_c[11] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1 ));
    NOR3C \scalestate_0/timecount_ret_58_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[0]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_130  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_94_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_142_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_130_Y ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_68_i ));
    OA1A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_6  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[3]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3_0 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_7 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[2]  (.A(
        \top_code_0_dumpdata_0[2] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[2] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_16  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[1] ), .C(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .Y(
        \timer_top_0/timer_0/N_17 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m34  
        (.A(\s_acq_change_0_s_stripnum[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[11]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i22_mux )
        );
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_60_i ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[9]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[8] ), 
        .Y(\DDS_0/dds_state_0/N_286 ));
    DFN1E1 \scalestate_0/CUTTIME90[5]  (.D(\top_code_0_scaledatain[5] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[5]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[9]  (.D(
        \DUMP_0/dump_coder_0/para4_4[9]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[9]_net_1 ));
    NOR3C \syn_md_module_1/syn_md_combine_0/syn_md_temp  (.A(
        scalestate_0_sw_acq1), .B(scalestate_0_rt_sw), .C(
        \syn_md_module_1/syn_md_combine_0/syn_md_temp_0_net_1 ), .Y(
        syn_md_tmp_c));
    DFN1 \state1ms_choice_0/reset_out  (.D(
        \state1ms_choice_0/reset_out_RNO_0_net_1 ), .CLK(GLA_net_1), 
        .Q(state1ms_choice_0_reset_out));
    NOR2A \DUMP_0/dump_state_0/cs_RNO_0[4]  (.A(
        \DUMP_0/dump_state_0/N_173 ), .B(
        \DUMP_0/dump_state_0/cs[3]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_185 ));
    AO1C \plusestate_0/CS_RNO_0[9]  (.A(\plusestate_0/CS[4]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst), .Y(
        \plusestate_0/CS_srsts_i_0[9] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[0]_net_1 ));
    DFN1 \DUMP_0/dump_coder_0/i[6]  (.D(
        \DUMP_0/dump_coder_0/i_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i[6] ));
    DFN1E1 \top_code_0/sd_sacq_data[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[5] ));
    NOR2B \scalestate_0/timecount_ret_66_RNO_0  (.A(
        \scalestate_0/CUTTIME180[14]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[14] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[4]  (.A(
        \scalestate_0/ACQ180_NUM[4]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[4]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_452 ));
    MX2B \plusestate_0/timecount_1_RNO[8]  (.A(\plusestate_0/N_79 ), 
        .B(\plusestate_0/N_215 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[8] ));
    DFN1E1 \top_code_0/sd_sacq_data[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[12] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[2]  (.D(
        \top_code_0_state_1ms_data[2] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[2]_net_1 ));
    MX2 \scalestate_0/load_out_RNO_0  (.A(\scalestate_0/N_1266 ), .B(
        scalestate_0_load_out), .S(\scalestate_0/N_1165 ), .Y(
        \scalestate_0/N_572 ));
    DFN1 \scalestate_0/CS[1]  (.D(\scalestate_0/CS_RNO_1[1] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[1]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[12]  (.A(
        \DDS_0/dds_state_0/para[12]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_329 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[12] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_3  (.A(
        \timer_top_0/timer_0/timedata[14]_net_1 ), .B(
        \timer_top_0/dataout[14] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_3_Y ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i22_mux ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datathree  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_1_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/un2_datathree ));
    AO1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_61  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_58_i ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_5_0 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_10_0 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[14]_net_1 ));
    NOR3C \top_code_0/k1_RNO_1  (.A(
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_4 ), .B(
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_3 ), .C(
        \top_code_0/N_11_3 ), .Y(\top_code_0/N_11 ));
    AO1A \scalestate_0/timecount_20_iv_5_RNO[11]  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[11]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[11] ), .Y(
        \scalestate_0/timecount_20_iv_0[11] ));
    AO1C \scalestate_0/necount_cmp_1/AO1C_0  (.A(
        \scalestate_0/necount[1]_net_1 ), .B(
        \scalestate_0/NE_NUM[1]_net_1 ), .C(
        \scalestate_0/necount[0]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/AO1C_0_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_149  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_75_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_127_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_149_Y ));
    NOR3C \scalestate_0/timecount_ret_67_RNO_1  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[14]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[14] ));
    OA1B \plusestate_0/CS_RNO[1]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[1]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[1] )
        , .Y(\plusestate_0/CS_RNO_0[1]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[5]  (.A(
        \DDS_0/dds_state_0/para[5]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_319 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[5] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m277  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_276 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_277 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_278 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[3]  (.A(
        \ClockManagement_0/long_timer_0/count_c2 ), .B(
        \ClockManagement_0/long_timer_0/count[3]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n3 ));
    AO1 \PLUSE_0/qq_state_1/Q1Q8_Q2Q7_RNO_0  (.A(\PLUSE_0/i_2[3] ), .B(
        \PLUSE_0/qq_state_1/cs[3]_net_1 ), .C(
        \PLUSE_0/qq_state_1/cs[4]_net_1 ), .Y(
        \PLUSE_0/qq_state_1/stateover_0_sqmuxa_i_0 ));
    DFN1 \s_acq_change_0/s_stripnum[3]  (.D(
        \s_acq_change_0/s_stripnum_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[3] ));
    IOIN_IB \ADC_pad[1]/U0/U1  (.YIN(\ADC_pad[1]/U0/NET1 ), .Y(
        \ADC_c[1] ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_51  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[7] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[8] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[10] )
        );
    IOPAD_IN \ADC_pad[4]/U0/U0  (.PAD(ADC[4]), .Y(\ADC_pad[4]/U0/NET1 )
        );
    MX2 \topctrlchange_0/soft_dump_RNO_0  (.A(soft_dump_net_0), .B(
        \topctrlchange_0/soft_dump_6 ), .S(\dds_change_0.un1_change_2 )
        , .Y(\topctrlchange_0/N_11 ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_0_i_i )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_8_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7_net_1 )
        );
    NOR2B \state_1ms_0/timecount_RNO_3[8]  (.A(
        \state_1ms_0/CUTTIME[8]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[8] ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_5  (.A(\ADC_c[5] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_5 ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_14  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] )
        , .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_5 ));
    DFN1 \DUMP_ON_0/off_on_timer_0/count[1]  (.D(
        \DUMP_ON_0/off_on_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/count_5[1] ));
    OA1B \top_code_0/pluseload_RNO_0  (.A(\top_code_0/N_161 ), .B(
        \top_code_0/N_175 ), .C(top_code_0_pluseload), .Y(
        \top_code_0/N_297 ));
    IOIN_IB \ADC_pad[11]/U0/U1  (.YIN(\ADC_pad[11]/U0/NET1 ), .Y(
        \ADC_c[11] ));
    DFN1E1 \top_code_0/dump_cho[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/dump_cho_1_sqmuxa ), .Q(
        \top_code_0_dump_cho_0[0] ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_41  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[3]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[8] ));
    NOR2A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[9]  (.A(
        \pd_pluse_top_0/i_0[5] ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_178 ));
    DFN1E1 \scanstate_0/acqtime[2]  (.D(\top_code_0_scandata[2] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[2]_net_1 ));
    OR3 \scalestate_0/timecount_20_iv_8[5]  (.A(
        \scalestate_0/timecount_20_iv_0[5] ), .B(
        \scalestate_0/OPENTIME_TEL_m[5] ), .C(
        \scalestate_0/timecount_20_iv_4[5]_net_1 ), .Y(
        \scalestate_0/timecount_20_iv_8[5]_net_1 ));
    XA1C \PLUSE_0/qq_coder_1/i_RNO_4[1]  (.A(\PLUSE_0/count_7[3] ), .B(
        \PLUSE_0/qq_para1[3] ), .C(\PLUSE_0/count_7[4] ), .Y(
        \PLUSE_0/qq_coder_1/i_0_0[1] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[3] ));
    DFN1E1 \plusestate_0/DUMPTIME[10]  (.D(\top_code_0_plusedata[10] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[10]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[19]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[19]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[19] ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/count_RNIV293[1]  (.A(
        \DSTimer_0/dump_sustain_timer_0/count[1]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_c1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m37  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_38_i ));
    IOPAD_TRI \relay_close_pad[5]/U0/U0  (.D(
        \relay_close_pad[5]/U0/NET1 ), .E(\relay_close_pad[5]/U0/NET2 )
        , .PAD(relay_close[5]));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i4_mux ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[1]  (.D(
        \top_code_0_pd_pluse_data[1] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[1]_net_1 ));
    IOPAD_IN \ADC_pad[8]/U0/U0  (.PAD(ADC[8]), .Y(\ADC_pad[8]/U0/NET1 )
        );
    OA1C \top_code_0/pd_pluse_load_RNO  (.A(\top_code_0/N_203 ), .B(
        top_code_0_pd_pluse_load), .C(\top_code_0/N_290 ), .Y(
        \top_code_0/N_82 ));
    DFN1 \timer_top_0/state_switch_0/clk_en_scale_0  (.D(
        \timer_top_0/state_switch_0/clk_en_scale_0_0_a6_0_a5_net_1 ), 
        .CLK(GLA_net_1), .Q(timer_top_0_clk_en_scale_0));
    NOR3 \DDS_0/dds_state_0/para_RNO[19]  (.A(
        \DDS_0/dds_state_0/N_508 ), .B(\DDS_0/dds_state_0/N_507 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[19] ), .Y(
        \DDS_0/dds_state_0/N_165 ));
    DFN1 \DUMP_ON_0/off_on_coder_0/i[0]  (.D(
        \DUMP_ON_0/off_on_coder_0/i_RNO_5[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/i_5[0] ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNIUJ9A[10]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[10]_net_1 ), .B(
        \sd_acq_top_0/i_0[8] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_233 ));
    DFN1E1 \scalestate_0/CUTTIME180[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[5]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_66_i ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[10]  (.D(
        \top_code_0_dds_configdata[9] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[10]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_9  (.A(\ADC_c[1] ), 
        .B(top_code_0_n_s_ctrl), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIGCUL3[2]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_5[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_4[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_11[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_13[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI0Q1G[6]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[6]_net_1 ), 
        .B(\pd_pluse_top_0/count_1[6] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_6[0] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[27]  (.A(
        \top_code_0_dds_configdata[10] ), .B(\DDS_0/dds_state_0/N_569 )
        , .C(\DDS_0/dds_state_0/N_474 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[27] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[4]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[4] ), 
        .CLK(GLA_net_1), .E(top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[4]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[7]  (.D(
        \top_code_0_pd_pluse_data[7] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[7]_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_12[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_11[4] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_13[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_15[4] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[25]  (.D(
        \top_code_0_dds_configdata[8] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[25]_net_1 ));
    AO1A \top_code_0/state_1ms_start_ret_3_RNO  (.A(\top_code_0/N_192 )
        , .B(\top_code_0/N_334 ), .C(\top_code_0/N_162 ), .Y(
        \top_code_0/N_112 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNILH9A4[9]  (.A(
        \ClockManagement_0/long_timer_0/count_c8 ), .B(
        \ClockManagement_0/long_timer_0/count[9]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c9 ));
    IOPAD_IN \xa_pad[9]/U0/U0  (.PAD(xa[9]), .Y(\xa_pad[9]/U0/NET1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[2] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_68_i ));
    OR3 \CAL_0/cal_div_0/count_RNIE3RN3[1]  (.A(
        \CAL_0/cal_div_0/clear_n4_NE_1 ), .B(
        \CAL_0/cal_div_0/clear_n4_NE_0 ), .C(
        \CAL_0/cal_div_0/clear_n4_NE_2 ), .Y(\CAL_0/cal_div_0/clear_n )
        );
    NOR2B \DUMP_0/dump_timer_0/count_RNO_1[11]  (.A(\DUMP_0/count[10] )
        , .B(\DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_23_0 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[7] ));
    DFN1E1 \top_code_0/s_addchoice_0[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_0[1] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[18]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[18]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_3[13]  (.A(
        \state_1ms_0/CUTTIME[13]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[13] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[11] ));
    DFN1E1 \scalestate_0/DUMPTIME[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[13]_net_1 ));
    NOR3A \DUMP_0/dump_coder_0/para19  (.A(\top_code_0_dump_cho_0[2] ), 
        .B(\top_code_0_dump_cho_0[0] ), .C(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para19_net_1 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[6]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c4 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n6 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_10_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ), .B(
        \sd_acq_top_0/count_1[9] ), .C(\sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_14_net ));
    DFN1E1 \noisestate_0/timecount_1[5]  (.D(
        \noisestate_0/timecount_5[5] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[5] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[31]  (.A(
        \DDS_0/dds_state_0/para_reg[31]_net_1 ), .B(
        \DDS_0/dds_state_0/N_535_0 ), .C(\DDS_0/dds_state_0/N_520 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_0[31] ));
    OR3A \top_code_0/sd_sacq_load_RNO_0  (.A(\xa_c[1] ), .B(
        \top_code_0/N_148 ), .C(\top_code_0/N_163 ), .Y(
        \top_code_0/N_195 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[4]_net_1 ));
    NOR2B \DUMP_0/dump_timer_0/count_RNO[10]  (.A(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_0/dump_timer_0/count_n10_tz ), .Y(
        \DUMP_0/dump_timer_0/count_n10 ));
    AOI1 \state_1ms_0/CS_i_RNO[0]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[9]_net_1 ), .C(\state_1ms_0/N_204s_i_i_0 ), .Y(
        \state_1ms_0/CS_i_RNO_1[0] ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m42_0 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[1]_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[30]  (.D(
        \top_code_0_dds_configdata[13] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[30]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m27  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_28 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_2_i ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[7]  (.A(
        \state_1ms_0_timecount[7] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_207 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m114  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[3] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_115 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[12]  (.D(
        \ClockManagement_0/long_timer_0/count_n12 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[12]_net_1 ));
    OR3C \CAL_0/cal_div_0/count_RNO[0]  (.A(net_33), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(
        \CAL_0/cal_div_0/count[0]_net_1 ), .Y(
        \CAL_0/cal_div_0/count_5[0] ));
    OR2A \scalestate_0/pn_out_RNO_1  (.A(\scalestate_0/N_1201 ), .B(
        top_code_0_pn_change), .Y(\scalestate_0/pn_out_4 ));
    NOR3C \timer_top_0/state_switch_0/clk_en_scan_RNO  (.A(net_27), .B(
        \timer_top_0/timer_0_time_up ), .C(top_code_0_scan_start), .Y(
        \timer_top_0/state_switch_0/clk_en_scan_RNO_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[9]  (.D(
        \DUMP_0/dump_coder_0/para2_4[9]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[9]_net_1 ));
    DFN1E1 \top_code_0/state_1ms_data[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[2] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m96  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_93 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_96 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_97 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs_i[0]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .CLK(ddsclkout_c), .Q(
        \pd_pluse_top_0/pd_pluse_state_0/cs_i[0]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_17  (.A(
        \timer_top_0/timer_0/N_17 ), .B(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .Y(
        \timer_top_0/timer_0/I_17_0 ));
    DFN1 \DUMP_0/dump_coder_0/i[3]  (.D(
        \DUMP_0/dump_coder_0/i_RNO_0[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_0[3] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[4]  (.A(
        \top_code_0_s_acqnum_2[4] ), .B(\scalestate_0_s_acqnum[4] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[4] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[12]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c10 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n12 ));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[3]  (.D(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[3] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/i_1[3] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIEAD6C[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_17[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_16[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_18[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE[0] ));
    DFN1 \scalestate_0/s_acqnum_1[3]  (.D(
        \scalestate_0/s_acqnum_1_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[3] ));
    DFN1 \s_acq_change_0/s_acqnum[7]  (.D(
        \s_acq_change_0/s_acqnum_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[7] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/dataout[12]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[12] ), .B(
        top_code_0_n_s_ctrl_1), .Y(\Signal_Noise_Acq_0_dataout[12] ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[6]  (.D(
        \top_code_0_state_1ms_data[6] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[6]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIQIEH[12]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[12]_net_1 )
        , .B(\pd_pluse_top_0/count[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_12[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIVMUE[6]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[6]_net_1 ), 
        .B(\pd_pluse_top_0/count_1[6] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_6[0] ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIB62L[10]  (.A(
        \DUMP_0/dump_coder_0/para4[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_10[0] ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIKQMS2[7]  (.A(
        \DUMP_0/dump_timer_0/count_c6 ), .B(\DUMP_0/count_0[7] ), .Y(
        \DUMP_0/dump_timer_0/count_c7 ));
    MX2 \noisestate_0/timecount_1_RNO[7]  (.A(\noisestate_0/N_64 ), .B(
        \noisestate_0/timecount_cnst[4] ), .S(\noisestate_0/N_228 ), 
        .Y(\noisestate_0/timecount_5[7] ));
    OA1A \DDS_0/dds_state_0/cs_RNO[5]  (.A(\DDS_0/dds_state_0/N_224 ), 
        .B(\DDS_0/dds_state_0/cs[4]_net_1 ), .C(
        \DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/cs_RNO[5]_net_1 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[2]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n2 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[7]  (.A(\scalestate_0/N_554 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[7]_net_1 ));
    NOR2A \ClockManagement_0/long_timer_0/count_RNO[0]  (.A(
        \ClockManagement_0/long_timer_0/en_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[0]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/N_95 ));
    AO1A \scalestate_0/timecount_ret_72_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[7]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[7] ), .Y(
        \scalestate_0/timecount_20_iv_1[7] ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_9  (.A(
        \scalestate_0/NE_NUM[4]_net_1 ), .B(
        \scalestate_0/necount[4]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_9_Y ));
    DFN1 \PLUSE_0/qq_timer_1/count[0]  (.D(
        \PLUSE_0/qq_timer_1/count_n0 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_7[0] ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_8  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_8_net_1 )
        );
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m31  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_32 ));
    NOR2B \scalestate_0/timecount_ret_54_RNO_0  (.A(
        \scalestate_0/CUTTIME180[19]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[19] ));
    OR2B \scalestate_0/long_opentime_RNO_1  (.A(
        \scalestate_0/CS[8]_net_1 ), .B(\scalestate_0/N_1196 ), .Y(
        \scalestate_0/N_1163 ));
    DFN1E1 \top_code_0/s_load  (.D(\top_code_0/N_94 ), .CLK(GLA_net_1), 
        .E(net_27), .Q(top_code_0_s_load));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_23  (.A(
        \timer_top_0/timer_0/N_15 ), .B(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .Y(
        \timer_top_0/timer_0/I_23_0 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m83  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_84 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[2]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_12_i ), .CLK(
        GLA_net_1), .E(top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[2]_net_1 ));
    IOPAD_TRI \syn_md_out_pad/U0/U0  (.D(\syn_md_out_pad/U0/NET1 ), .E(
        \syn_md_out_pad/U0/NET2 ), .PAD(syn_md_out));
    AO1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[12]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .B(
        \sd_acq_top_0/i[9] ), .C(\sd_acq_top_0/sd_sacq_state_0/cs4 ), 
        .Y(\sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[12] ));
    DFN1 \scalestate_0/strippluse[8]  (.D(
        \scalestate_0/strippluse_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[8] ));
    NOR3C \PLUSE_0/bri_timer_0/count_RNIM4N5[0]  (.A(
        \PLUSE_0/count_8[1] ), .B(\PLUSE_0/count_8[0] ), .C(
        \PLUSE_0/count_8[2] ), .Y(\PLUSE_0/bri_timer_0/count_c2 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIQ77S[11]  (
        .A(\pd_pluse_top_0/count_0[11] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[11]_net_1 ), 
        .C(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_8[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_1[0] ));
    DFN1 \DUMP_0/dump_timer_0/count[0]  (.D(
        \DUMP_0/dump_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_1[0] ));
    OR3 \scalestate_0/timecount_RNO[21]  (.A(
        \scalestate_0/timecount_20_0_iv_0[21] ), .B(
        \scalestate_0/OPENTIME_TEL_m[21] ), .C(
        \scalestate_0/timecount_20_0_iv_1[21] ), .Y(
        \scalestate_0/timecount_20[21] ));
    NOR2B \DDS_0/dds_state_0/para_RNO_0[35]  (.A(
        \DDS_0/dds_state_0/para[36]_net_1 ), .B(
        \DDS_0/dds_state_0/N_534 ), .Y(\DDS_0/dds_state_0/N_526 ));
    OR2B \DUMP_0/off_on_state_0/state_over_RNO  (.A(
        \DUMP_0/off_on_state_0/N_12_mux ), .B(
        state1ms_choice_0_reset_out), .Y(\DUMP_0/off_on_state_0/N_9 ));
    OR3 \top_code_0/plusedata_1_sqmuxa_0_o2_0  (.A(\xa_c[6] ), .B(
        \top_code_0/N_137 ), .C(\xa_c[5] ), .Y(\top_code_0/N_139 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[6]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_17_0 ), .Y(
        \timer_top_0/timer_0/timedata_4[6] ));
    NOR2 \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[5]  (.A(\i_6[1] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_217 ));
    NOR3C \scalestate_0/timecount_ret_72_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[7]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[7] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m275  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_276 ));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[4]  (.D(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[4]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/i_0[4] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[8]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[8] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_0[8] ));
    OR3A \top_code_0/pluse_noise_ctrl_3_i_o2  (.A(\xa_c[7] ), .B(
        \top_code_0/N_139 ), .C(\top_code_0/N_154 ), .Y(
        \top_code_0/N_176 ));
    AO1 \scalestate_0/timecount_ret_59_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[0]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[0] ), .Y(
        \scalestate_0/timecount_20_iv_4[0] ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_70_i ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNIOS8L2[8]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c6 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c8 ));
    AO1C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_17  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_2 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_8 ));
    DFN1E1 \scalestate_0/timecount_ret_33  (.D(
        \scalestate_0/timecount_m1_e_2_2 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_m1_e_2_2_reto ));
    DFN1 \noisestate_0/soft_d  (.D(\noisestate_0/soft_d_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(noisestate_0_soft_d));
    MX2 \scanstate_0/timecount_1_RNO_0[7]  (.A(
        \scanstate_0/acqtime[7]_net_1 ), .B(
        \scanstate_0/dectime[7]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_65 ));
    DFN1E1 \noisestate_0/acqtime[9]  (.D(\top_code_0_noisedata[9] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[9]_net_1 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[0]  (.A(
        \top_code_0_dumpdata_0[0] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[0] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[3]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[3] ));
    NOR3C \DDS_0/dds_coder_0/i_RNO[2]  (.A(
        \DDS_0/dds_coder_0/N_18_mux ), .B(
        \DDS_0/dds_coder_0/m12_2_net_1 ), .C(\DDS_0/count[2] ), .Y(
        \DDS_0/dds_coder_0/i_RNO[2]_net_1 ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_0  (.A(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .B(
        \timer_top_0/dataout[21] ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR2A_0_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_0_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIFU6T[19]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[19]_net_1 ), .B(
        \sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_19[0] ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/NE_NUM[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_3_Y ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[10]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[10] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[10]_net_1 ));
    DFN1 \top_code_0/state_1ms_start_ret_2  (.D(\top_code_0/un1_xa_4 ), 
        .CLK(GLA_net_1), .Q(\top_code_0/un1_xa_4_reto ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_61  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[28] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[13] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[15] ), .Y(
        \timer_top_0/timer_0/N_2 ));
    DFN1E1 \scalestate_0/DUMPTIME[4]  (.D(\top_code_0_scaledatain[4] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[4]_net_1 ));
    NOR2A \PLUSE_0/bri_state_0/cs_RNO_10[3]  (.A(
        \PLUSE_0/bri_state_0/cs[1]_net_1 ), .B(\PLUSE_0/i_3[2] ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_1_0 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[6]_net_1 ));
    DFN1E1 \top_code_0/state_1ms_data[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[15] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[1]  (.A(
        \noisestate_0_timecount[1] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_235 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_60_i ));
    NOR2B \scalestate_0/timecount_ret_49_RNO  (.A(
        \scalestate_0/OPENTIME_TEL[17]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[17] ));
    DFN1 \syn_md_module_1/syn_md_0/syn_md_out  (.D(
        \syn_md_module_1/syn_md_0/N_14 ), .CLK(GLA_net_1), .Q(
        syn_md_out_c));
    MX2 \state_1ms_0/timecount_RNO_0[19]  (.A(
        \state_1ms_0/timecount_8[19] ), .B(\state_1ms_0_timecount[19] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_86 ));
    DFN1E1 \state_1ms_0/PLUSETIME[8]  (.D(
        \top_code_0_state_1ms_data[8] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[8]_net_1 ));
    AND2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/VAND2_17_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_24_net ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNI3RUE[8]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[8]_net_1 ), 
        .B(\pd_pluse_top_0/count_0[8] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_8[0] ));
    DFN1E1 \top_code_0/dumpload  (.D(\top_code_0/N_70 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_dumpload));
    DFN1 \scalestate_0/strippluse[9]  (.D(
        \scalestate_0/strippluse_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[9] ));
    OR3 \DUMP_0/dump_state_0/cs_RNO_2[5]  (.A(
        \DUMP_0/dump_state_0/N_201 ), .B(
        \DUMP_0/dump_state_0/cs[6]_net_1 ), .C(
        \DUMP_0/dump_state_0/N_203 ), .Y(\DUMP_0/dump_state_0/N_167 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_6 ), .B(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_1_sqmuxa ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_41 ));
    AO1 \state_1ms_0/timecount_RNO_4[14]  (.A(
        \state_1ms_0/S_DUMPTIME[14]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[14] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[14] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_60_i ));
    NOR3B \scalestate_0/timecount_ret_27_RNO  (.A(
        \scalestate_0/timecount_11_sqmuxa ), .B(\scalestate_0/N_1089 ), 
        .C(\scalestate_0/N_258_0 ), .Y(\scalestate_0/timecount_m3_e_1 )
        );
    NOR2B \ClockManagement_0/long_timer_0/count_RNI02OQ4[8]  (.A(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_7 ), .B(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_6 ), .Y(
        \ClockManagement_0/long_timer_0/count_c11 ));
    DFN1 \PLUSE_0/qq_state_1/cs[2]  (.D(
        \PLUSE_0/qq_state_1/cs_RNO_2[2] ), .CLK(GLA_net_1), .Q(Q4Q5_c));
    NOR2B \scalestate_0/necount_RNO[9]  (.A(\scalestate_0/N_739 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[9]_net_1 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[5]  (.D(
        \top_code_0_state_1ms_data[5] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[5]_net_1 ));
    XO1 \PLUSE_0/qq_coder_1/i_reg10_NE_2[0]  (.A(\PLUSE_0/count_7[1] ), 
        .B(\PLUSE_0/qq_para3[1] ), .C(
        \PLUSE_0/qq_coder_1/i_reg10_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_NE_2[0]_net_1 ));
    DFN1E1 \noisestate_0/timecount_1[2]  (.D(
        \noisestate_0/timecount_5[2] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[2] ));
    NOR2B \DUMP_OFF_1/off_on_timer_0/count_RNISQ1I[2]  (.A(
        \DUMP_OFF_1/off_on_timer_0/count_c1 ), .B(
        \DUMP_OFF_1/count_4[2] ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_c2 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[10]  (.A(
        \s_acq_change_0/N_66 ), .B(net_27), .Y(
        \s_acq_change_0/s_stripnum_RNO[10]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[13]_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[3]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[3] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[3] ));
    DFN1E1 \top_code_0/scaledatain[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[10] ));
    OA1B \plusestate_0/CS_RNO[5]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[5]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[5] )
        , .Y(\plusestate_0/CS_RNO_0[5]_net_1 ));
    NOR3C \scalestate_0/STRIPNUM90_NUM_1_sqmuxa_0_a2  (.A(
        \top_code_0_scalechoice_0_0[0] ), .B(\scalestate_0/N_60 ), .C(
        \scalestate_0/N_67 ), .Y(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[7]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[7] ));
    DFN1 \PLUSE_0/qq_coder_1/i[0]  (.D(\PLUSE_0/qq_coder_1/i_RNO_8[0] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_7[0] ));
    OR2A \scalestate_0/CS_RNI62781[17]  (.A(\scalestate_0/N_1194 ), .B(
        \scalestate_0/N_1265 ), .Y(\scalestate_0/N_1209 ));
    OA1C \top_code_0/scaleload_RNO  (.A(\top_code_0/N_217 ), .B(
        top_code_0_scaleload), .C(\top_code_0/N_304 ), .Y(
        \top_code_0/N_96 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIS1KD[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_4[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_3[0] ));
    DFN1 \n_acq_change_0/n_acq_start  (.D(
        \n_acq_change_0/n_acq_start_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        n_acq_change_0_n_acq_start));
    OR3 \scalestate_0/timecount_ret_85_RNO  (.A(
        \scalestate_0/PLUSETIME90_m[11] ), .B(
        \scalestate_0/DUMPTIME_m[11] ), .C(
        \scalestate_0/S_DUMPTIME_m[11] ), .Y(
        \scalestate_0/timecount_20_iv_6[11] ));
    DFN1 \DUMP_0/dump_state_0/off_start  (.D(
        \DUMP_0/dump_state_0/off_start_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(\DUMP_0/dump_state_0_off_start ));
    NOR2B \state1ms_choice_0/pluse_start_RNO  (.A(
        \state1ms_choice_0/pluse_start_5 ), .B(net_27), .Y(
        \state1ms_choice_0/pluse_start_RNO_1 ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[5]  (.A(
        \top_code_0_dumpdata_0[5] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[5]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO[11]  (.A(\state_1ms_0/N_78 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[11]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m247  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_246 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_247 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_248 ));
    NOR2A \top_code_0/dds_configdata_1_sqmuxa_0_a2_1  (.A(net_27), .B(
        \top_code_0/N_147 ), .Y(\top_code_0/dds_configdata_1_sqmuxa_1 )
        );
    NOR2A \noisestate_0/acqtime_1_sqmuxa  (.A(top_code_0_nstateload), 
        .B(top_code_0_nstatechoice), .Y(
        \noisestate_0/acqtime_1_sqmuxa_net_1 ));
    DFN1 \state_1ms_0/timecount[6]  (.D(
        \state_1ms_0/timecount_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[6] ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_24  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_46_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[0] )
        );
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[11]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n11 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ));
    OR2A \scanstate_0/CS_RNIMKVU[6]  (.A(net_33), .B(
        \scanstate_0/N_255 ), .Y(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ));
    NOR2B \state_1ms_0/timecount_RNO[13]  (.A(\state_1ms_0/N_80 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[13]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[18]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[18]_net_1 ));
    NOR2B \nsctrl_choice_0/dumpon_ctr_RNO  (.A(
        \nsctrl_choice_0/dumpon_ctr_5 ), .B(net_27), .Y(
        \nsctrl_choice_0/dumpon_ctr_RNO_0_net_1 ));
    DFN1E1 \scanstate_0/timecount_1[13]  (.D(
        \scanstate_0/timecount_5[13] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[13] ));
    IOBI_IB_OB_EB \xd_pad[4]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[4] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[4]/U0/NET3 ), .DOUT(\xd_pad[4]/U0/NET1 ), .EOUT(
        \xd_pad[4]/U0/NET2 ), .Y(\xd_in[4] ));
    DFN1 \timer_top_0/timer_0/timedata[17]  (.D(
        \timer_top_0/timer_0/timedata_4[17] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[17]_net_1 ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y ));
    AO1C \DUMP_0/dump_state_0/timer_start_RNO_1  (.A(\DUMP_0/i_2[1] ), 
        .B(\DUMP_0/dump_state_0/cs[3]_net_1 ), .C(
        \DUMP_0/dump_state_0/N_173 ), .Y(\DUMP_0/dump_state_0/ns[3] ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[2]  (.A(
        \s_acq_change_0/s_stripnum_5[2] ), .B(
        \s_acq_change_0_s_stripnum[2] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_58 ));
    AO1 \state_1ms_0/timecount_RNO_4[12]  (.A(
        \state_1ms_0/S_DUMPTIME[12]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[12] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[12] ));
    NOR2A \PLUSE_0/qq_timer_0/count_RNO[0]  (.A(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ), .B(
        \PLUSE_0/count_9[0] ), .Y(\PLUSE_0/qq_timer_0/count_n0 ));
    NOR3C \top_code_0/un1_state_1ms_rst_n117_43_i_a2_1_1  (.A(
        \xa_c[2] ), .B(\top_code_0/N_329 ), .C(\xa_c[4] ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_43_i_a2_1_1_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m64  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_61 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_64 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_65 ));
    OR3B \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[12]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .B(
        \sd_acq_top_0/i_5[3] ), .C(\sd_acq_top_0/i_5[2] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_208 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m42_1 ));
    DFN1E1 \noisestate_0/acqtime[6]  (.D(\top_code_0_noisedata[6] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[6]_net_1 ));
    IOPAD_IN \ADC_pad[5]/U0/U0  (.PAD(ADC[5]), .Y(\ADC_pad[5]/U0/NET1 )
        );
    NOR2B \top_code_0/k2_RNO  (.A(\top_code_0/N_806 ), .B(net_27), .Y(
        \top_code_0/k2_RNO_net_1 ));
    DFN1E1 \state_1ms_0/CUTTIME[5]  (.D(\top_code_0_state_1ms_data[5] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[5]_net_1 ));
    OA1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[2]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[2]_net_1 ), .B(
        \sd_acq_top_0/i_2[4] ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs[1]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_214 ));
    NOR2 \sd_acq_top_0/sd_sacq_state_0/cs_RNIH512[14]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[14]_net_1 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[15]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/ns_0_1_i_a2_0 ));
    DFN1 \scalestate_0/s_acqnum_1[1]  (.D(
        \scalestate_0/s_acqnum_1_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[1] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIC2DM[1]  (.A(
        \sd_acq_top_0/count_10[1] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[1]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_9[0] ));
    AND2 \ClockManagement_0/clk_10k_0/un1_count_1_I_53  (.A(
        \ClockManagement_0/clk_10k_0/count[4]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_1[0] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[3]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[3] ));
    DFN1 \noisestate_0/dumpoff_ctr  (.D(
        \noisestate_0/dumpoff_ctr_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        noisestate_0_dumpoff_ctr));
    NOR2B \DUMP_0/dump_state_0/cs_RNO[1]  (.A(
        \DUMP_0/dump_state_0/N_171 ), .B(\DUMP_0/dump_state_0/cs4 ), 
        .Y(\DUMP_0/dump_state_0/cs_nsss[1] ));
    NOR2B \bridge_div_0/clk_4f_reg2_RNIREDC  (.A(
        \bridge_div_0/clk_4f_reg1_net_1 ), .B(
        \bridge_div_0/clk_4f_reg2_i_0 ), .Y(clk_4f_en));
    NOR2B \top_code_0/inv_turn_RNO  (.A(\top_code_0/N_802 ), .B(net_27)
        , .Y(\top_code_0/inv_turn_RNO_net_1 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/YAND2_22_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_16_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net ), 
        .C(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_27_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_18  
        (.A(\s_acq_change_0_s_stripnum[3] ), .B(
        \s_acq_change_0_s_stripnum[4] ), .C(
        \s_acq_change_0_s_stripnum[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] )
        );
    XOR2 \DUMP_0/dump_coder_0/para5_RNIEC8P[11]  (.A(
        \DUMP_0/dump_coder_0/para5[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_11[0] ));
    NOR3C \DUMP_0/dump_state_0/cs_RNIM9N51[6]  (.A(
        \DUMP_0/dump_state_0/N_166 ), .B(\DUMP_0/dump_state_0/N_206 ), 
        .C(\DUMP_0/dump_state_0/cs4 ), .Y(
        \DUMP_0/dump_state_0/cs_nsss[6] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m53  
        (.A(\s_acq_change_0_s_stripnum[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[5]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i8_mux ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_54_i ));
    DFN1E1 \top_code_0/scanload  (.D(\top_code_0/N_100 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_scanload));
    OR3 \scalestate_0/timecount_ret_56_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[19] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[19] ), .C(
        \scalestate_0/timecount_20_0_iv_2[19] ), .Y(
        \scalestate_0/timecount_20_0_iv_4[19] ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_11  (.A(
        \scalestate_0/NE_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_5 ));
    MX2 \PLUSE_0/bri_state_0/up/U0  (.A(\PLUSE_0/up ), .B(
        \PLUSE_0/bri_state_0/down30 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/up/Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[6]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[6]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_276 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[8]  (.A(
        \noisestate_0_timecount[8] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_245 ));
    OA1C \top_code_0/bridge_load_0_RNIBM406  (.A(\top_code_0/N_216 ), 
        .B(top_code_0_bridge_load_0), .C(\top_code_0/N_270 ), .Y(
        \top_code_0/N_62 ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_8[10]  (.A(
        \sd_acq_top_0/count[20] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[20]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_17[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_1[10] ));
    AO1A \state_1ms_0/timecount_RNO_4[5]  (.A(
        \state_1ms_0/S_DUMPTIME[5]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CUTTIME_i_m[5] ), 
        .Y(\state_1ms_0/timecount_8_iv_2[5] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m41_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[18] ));
    AND3 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_1_7_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/count_1[6] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_7_net ));
    DFN1 \scalestate_0/CS[6]  (.D(\scalestate_0/CS_RNO_1[6] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[6]_net_1 ));
    NOR3 \DUMP_0/dump_coder_0/para15  (.A(\top_code_0_dump_cho_0[2] ), 
        .B(\top_code_0_dump_cho_0[0] ), .C(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para15_net_1 ));
    IOPAD_BI \xd_pad[9]/U0/U0  (.D(\xd_pad[9]/U0/NET1 ), .E(
        \xd_pad[9]/U0/NET2 ), .Y(\xd_pad[9]/U0/NET3 ), .PAD(xd[9]));
    DFN1 \state_1ms_0/reset_out  (.D(\state_1ms_0/reset_out_RNO_1 ), 
        .CLK(GLA_net_1), .Q(state_1ms_0_reset_out));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[4]  (.D(
        \top_code_0_pd_pluse_data[4] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[4]_net_1 ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_10[10]  (.A(
        \sd_acq_top_0/count_3[6] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[6]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_4[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_8[10] ));
    NOR2B \DDS_0/dds_state_0/para_RNO_0[0]  (.A(
        \DDS_0/dds_state_0/para[1]_net_1 ), .B(
        \DDS_0/dds_state_0/N_534 ), .Y(\DDS_0/dds_state_0/N_528 ));
    DFN1 \scalestate_0/CS[18]  (.D(\scalestate_0/CS_RNO[18]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[18]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m85  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_84 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_85 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_86 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[5]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c4 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n5 ));
    DFN1C0 \bridge_div_0/clk_4f_reg1  (.D(\bridge_div_0/clk_4f ), .CLK(
        ddsclkout_c), .CLR(bri_dump_sw_0_reset_out_0), .Q(
        \bridge_div_0/clk_4f_reg1_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_164  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_164_Y ));
    MX2 \scalestate_0/CS_RNO_0[9]  (.A(\scalestate_0/CS[9]_net_1 ), .B(
        \scalestate_0/CS[8]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1223 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_16[3]  (.A(
        \DUMP_0/dump_coder_0/para1[6]_net_1 ), .B(\DUMP_0/count_0[6] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_6[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m46_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[13] ));
    OR3 \scalestate_0/timecount_ret_31_RNIC8I  (.A(
        \scalestate_0/timecount_20_iv_3_reto[4] ), .B(
        \scalestate_0/timecount_20_iv_2_reto[4] ), .C(
        \scalestate_0/timecount_20_iv_6_reto[4] ), .Y(
        \scalestate_0/timecount_20_iv_9_reto[4] ));
    AND2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y ));
    OR2A \PLUSE_0/bri_state_0/csse_10_0_o2  (.A(\PLUSE_0/i_3[2] ), .B(
        \PLUSE_0/i_8[1] ), .Y(\PLUSE_0/bri_state_0/N_142 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_26[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_5[0] ));
    DFN1E1 \top_code_0/state_1ms_data[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[4] ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_9_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_11_net ), 
        .B(\pd_pluse_top_0/count_0[11] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[11] ));
    DFN1E1 \scalestate_0/timecount_ret_2  (.D(
        \scalestate_0/timecount_20_iv_9[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_9_reto[6] ));
    NOR3A \PLUSE_0/qq_state_0/cs_RNO[3]  (.A(\PLUSE_0/qq_state_0/cs4 ), 
        .B(\PLUSE_0/qq_state_0/N_86 ), .C(\PLUSE_0/qq_state_0/N_87 ), 
        .Y(\PLUSE_0/qq_state_0/cs_RNO_1[3]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_data[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[15] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m24  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_25 ));
    DFN1 \top_code_0/noise_start_ret  (.D(top_code_0_noise_start), 
        .CLK(GLA_net_1), .Q(\top_code_0/top_code_0_noise_start_reto ));
    DFN1E1 \top_code_0/dumpdata[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[0] ));
    DFN1E1 \top_code_0/sigtimedata[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[14] ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[14]  (.A(\s_acq_change_0/N_84 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[14]_net_1 ));
    DFN1 \state1ms_choice_0/bri_cycle  (.D(
        \state1ms_choice_0/bri_cycle_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        state1ms_choice_0_bri_cycle));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[6]  (.A(
        \top_code_0_s_acqnum_2[6] ), .B(\scalestate_0_s_acqnum[6] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[6] ));
    MX2 \bri_dump_sw_0/dumpoff_ctr_RNO_0  (.A(plusestate_0_tetw_pluse), 
        .B(scalestate_0_dumpoff_ctr), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/dumpoff_ctr_5 ));
    AO1 \state_1ms_0/timecount_RNO_2[7]  (.A(
        \state_1ms_0/M_DUMPTIME[7]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[7] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[7] ));
    OR2A \DDS_0/dds_state_0/cs_RNO_1[2]  (.A(
        \DDS_0/dds_state_0/cs[2]_net_1 ), .B(\DDS_0/i[2] ), .Y(
        \DDS_0/dds_state_0/N_225 ));
    NOR2 \GPMI_0/xwe_xzcs2_syn_0/code_en_RNO_0  (.A(zcs2_c), .B(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_net_1 ), .Y(
        \GPMI_0/xwe_xzcs2_syn_0/code_en_0_0 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[0]  (.A(
        \top_code_0_s_acqnum_2[0] ), .B(\scalestate_0_s_acqnum[0] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[0] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[2] ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_7  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_0_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_6_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_16_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_7_Y ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNI9GII[0]  (.A(
        \DUMP_0/dump_coder_0/para4[0]_net_1 ), .B(\DUMP_0/count_1[0] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_0_0[0] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_8  (.A(\ADC_c[2] ), 
        .B(top_code_0_n_s_ctrl), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ));
    OA1B \state_1ms_0/CS_RNO[1]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[1]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[1] ), 
        .Y(\state_1ms_0/CS_RNO_3[1] ));
    AO1C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_5  (
        .A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[1]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_4_0 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_6 ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_26  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[4]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[0] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIAS6K[1]  (.A(
        \sd_acq_top_0/count_10[1] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[1]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_9[0] ));
    NOR2B \scalestate_0/timecount_ret_56_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[19]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[19] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[4] ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[5]  (.A(
        \ClockManagement_0/long_timer_0/count_c4 ), .B(
        \ClockManagement_0/long_timer_0/count[5]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n5 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[3]  (.A(\s_acq_change_0/N_59 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[3]_net_1 ));
    NOR3B \bridge_div_0/count_RNIHPOM7[3]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[3]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIHPOM7[3]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[3]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[3] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_11_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_11_net ));
    DFN1 \plusestate_0/CS[3]  (.D(\plusestate_0/CS_RNO_0[3]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[3]_net_1 ));
    IOPAD_TRI \relay_on_pad[1]/U0/U0  (.D(\relay_on_pad[1]/U0/NET1 ), 
        .E(\relay_on_pad[1]/U0/NET2 ), .PAD(relay_on[1]));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIDEET[10]  (.A(
        \DUMP_0/dump_coder_0/para6[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_10[0] ));
    MX2 \scalestate_0/CS_RNO_0[3]  (.A(\scalestate_0/CS[3]_net_1 ), .B(
        \scalestate_0/CS[2]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1218 ));
    NOR2B \scalestate_0/timecount_ret_57_RNO_1  (.A(
        \scalestate_0/OPENTIME[0]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[0] ));
    NOR3C \state_1ms_0/CUTTIME_161_e  (.A(\state_1ms_0/N_16 ), .B(
        \state_1ms_0/un1_PLUSECYCLE13_i_a2_0_net_1 ), .C(
        \top_code_0_state_1ms_lc[0] ), .Y(\state_1ms_0/N_380 ));
    NOR3A 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa_0_a2_0  
        (.A(top_code_0_pd_pluse_load), .B(
        \top_code_0_pd_pluse_choice[3] ), .C(
        \top_code_0_pd_pluse_choice[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/N_12 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m50  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_43 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_50 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_51 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_37_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_81  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_135_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_28_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_81_Y ));
    NOR3C \timer_top_0/state_switch_0/clk_en_noise_RNO  (.A(net_27), 
        .B(\timer_top_0/timer_0_time_up ), .C(top_code_0_noise_start), 
        .Y(\timer_top_0/state_switch_0/clk_en_noise_RNO_net_1 ));
    IOPAD_IN \OCX40MHz_pad/U0/U0  (.PAD(OCX40MHz), .Y(OCX40MHz_c));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_93  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_93_Y ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[5]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[5] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[5]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO[6]  (.A(\noisestate_0/N_63 ), .B(
        \noisestate_0/timecount_cnst[2] ), .S(\noisestate_0/N_228 ), 
        .Y(\noisestate_0/timecount_5[6] ));
    NOR2B \DDS_0/dds_state_0/para_reg_100_e  (.A(top_code_0_dds_choice)
        , .B(top_code_0_dds_load), .Y(\DDS_0/dds_state_0/N_569 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_1  (.A(\xd_in[13] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[13] ));
    DFN1 \state_1ms_0/CS[2]  (.D(\state_1ms_0/CS_RNO_3[2] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[2]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m245  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_246 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[9]_net_1 ));
    NOR3A \topctrlchange_0/interupt_RNO_4  (.A(
        nsctrl_choice_0_intertodsp), .B(\top_code_0_change_0[0] ), .C(
        \top_code_0_change_0[1] ), .Y(\topctrlchange_0/interin1_m ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_132  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_132_Y ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_7  (.A(\xd_in[7] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[7] ));
    DFN1 \state_1ms_0/timecount[15]  (.D(
        \state_1ms_0/timecount_RNO[15]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[15] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[16]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[16]_net_1 ));
    NOR2A \scalestate_0/fst_lst_pulse_RNI6R4S  (.A(
        \scalestate_0/N_297 ), .B(\scalestate_0/fst_lst_pulse_net_1 ), 
        .Y(\scalestate_0/sw_acq1_1_sqmuxa ));
    IOPAD_IN \ADC_pad[6]/U0/U0  (.PAD(ADC[6]), .Y(\ADC_pad[6]/U0/NET1 )
        );
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[2] ));
    NOR3C \scalestate_0/timecount_ret_11_RNO_1  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[7]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[7] ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[10]  (.A(\s_acq_change_0/N_80 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[10]_net_1 ));
    IOPAD_TRI \relay_close_pad[1]/U0/U0  (.D(
        \relay_close_pad[1]/U0/NET1 ), .E(\relay_close_pad[1]/U0/NET2 )
        , .PAD(relay_close[1]));
    DFN1E0 \DUMP_0/dump_coder_0/para3[1]  (.D(
        \DUMP_0/dump_coder_0/para4_4[1]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[1]_net_1 ));
    AX1C \scalestate_0/necount_inc_0/XOR2_2_1_inst  (.A(
        \scalestate_0/necount[0]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .C(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/necount1[2] ));
    OA1B \noisestate_0/CS_RNO[1]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[1]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[1] )
        , .Y(\noisestate_0/CS_RNO[1]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIUFCH[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[10]_net_1 ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_10[0] ));
    DFN1E1 \scalestate_0/CUTTIME180[19]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1661 ), .Q(\scalestate_0/CUTTIME180[19]_net_1 )
        );
    DFN1 \top_code_0/noise_rst  (.D(
        \top_code_0/noise_rst_0_0_RNIDOO43_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_noise_rst));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[12]  (.D(
        \top_code_0_pd_pluse_data[12] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[12]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[8]_net_1 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[9]  (.A(\scalestate_0/N_457 ), 
        .B(\scalestate_0/ACQECHO_NUM[9]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[9] ));
    DFN1E1 \scalestate_0/OPENTIME[1]  (.D(\top_code_0_scaledatain[1] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[1]_net_1 ));
    AOI1 \scalestate_0/necount_cmp_1/AOI1_ALEB  (.A(
        \scalestate_0/necount_cmp_1/AND3_0_Y ), .B(
        \scalestate_0/necount_cmp_1/AO1_1_Y ), .C(
        \scalestate_0/necount_cmp_1/AO1_0_Y ), .Y(
        \scalestate_0/necount_LE_NE_1 ));
    OR2B \noisestate_0/CS_RNIUO68[4]  (.A(\noisestate_0/CS[4]_net_1 ), 
        .B(top_code_0_noise_rst), .Y(\noisestate_0/N_191 ));
    OA1B \scanstate_0/CS_RNO[6]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[6]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[6] ), 
        .Y(\scanstate_0/CS_RNO_2[6] ));
    NOR2A \scanstate_0/acqtime_1_sqmuxa  (.A(top_code_0_scanload), .B(
        top_code_0_scanchoice), .Y(
        \scanstate_0/acqtime_1_sqmuxa_net_1 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_0  (.A(
        \timer_top_0/dataout[9] ), .B(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_0_Y ));
    IOIN_IB \XRD_pad/U0/U1  (.YIN(\XRD_pad/U0/NET1 ), .Y(XRD_c));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_39_i ));
    AND3B \DDS_0/dds_coder_0/m12_2  (.A(\DDS_0/count[6] ), .B(
        \DDS_0/count[5] ), .C(\DDS_0/dds_coder_0/m12_0_net_1 ), .Y(
        \DDS_0/dds_coder_0/m12_2_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m93  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_94 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/ADD_20x20_slow_I19_Y_1 )
        );
    MX2 \scalestate_0/s_acqnum_1_RNO_2[6]  (.A(
        \scalestate_0/ACQ180_NUM[6]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[6]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_454 ));
    AO1C \scalestate_0/dds_conf_RNO_1  (.A(\scalestate_0/un1_CS_20 ), 
        .B(\scalestate_0/N_1262 ), .C(timer_top_0_clk_en_scale), .Y(
        \scalestate_0/N_1173 ));
    DFN1E1 \bridge_div_0/dataall[2]  (.D(\bridge_div_0/dataall_1[2] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/dataall[2]_net_1 ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[0]  (.A(
        scalestate_0_s_acq), .B(net_27), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_9[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[2] ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/count[1]  (.D(
        \DSTimer_0/dump_sustain_timer_0/count_n1 ), .CLK(clock_10khz), 
        .Q(\DSTimer_0/dump_sustain_timer_0/count[1]_net_1 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_24  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[3] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[4] )
        );
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_6  (.A(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .B(
        \timer_top_0/dataout[16] ), .C(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_6_Y ));
    OR2A \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_RNO  (
        .A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_RNO_net_1 )
        );
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIAJEN[14]  (.A(
        \sd_acq_top_0/count_0[14] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[14]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_8[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_0[0] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[5]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n5 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ));
    XA1C \PLUSE_0/qq_coder_1/i_RNO_1[1]  (.A(\PLUSE_0/count_7[2] ), .B(
        \PLUSE_0/qq_para1[2] ), .C(\PLUSE_0/qq_coder_1/un1_count_1[0] )
        , .Y(\PLUSE_0/qq_coder_1/i_0_1[1] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[9]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c8 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n9 ));
    OAI1 \plusestate_0/timecount_1_RNO_1[4]  (.A(
        \plusestate_0/CS[8]_net_1 ), .B(\plusestate_0/CS[3]_net_1 ), 
        .C(top_code_0_pluse_rst_0), .Y(\plusestate_0/N_249 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i20_mux ));
    IOIN_IB \tri_ctrl_pad/U0/U1  (.YIN(\tri_ctrl_pad/U0/NET1 ), .Y(
        tri_ctrl_c));
    NOR2B \scalestate_0/necount_RNO[7]  (.A(\scalestate_0/N_737 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[7]_net_1 ));
    AO1 \scalestate_0/necount_cmp_1/AO1_1  (.A(
        \scalestate_0/necount_cmp_1/AND3_2_Y ), .B(
        \scalestate_0/necount_cmp_1/NAND3A_4_Y ), .C(
        \scalestate_0/necount_cmp_1/NAND3A_0_Y ), .Y(
        \scalestate_0/necount_cmp_1/AO1_1_Y ));
    INV \bridge_div_0/count_5_I_4  (.A(
        \bridge_div_0/count_RNIEMOM7[0]_net_1 ), .Y(
        \bridge_div_0/count_5[0] ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[8]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[8] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_8_inst ), .S(top_code_0_n_s_ctrl_1), 
        .Y(\Signal_Noise_Acq_0_dataout[8] ));
    DFN1 \DDS_0/dds_state_0/cs_i[0]  (.D(\DDS_0/dds_state_0/N_223 ), 
        .CLK(GLA_net_1), .Q(\DDS_0/dds_state_0/cs_i[0]_net_1 ));
    DFN1E1 \state_1ms_0/CUTTIME[8]  (.D(\top_code_0_state_1ms_data[8] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[8]_net_1 ));
    DFN1E1 \scalestate_0/DUMPTIME[1]  (.D(\top_code_0_scaledatain[1] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[1]_net_1 ));
    NOR3C \ClockManagement_0/long_timer_0/count_RNIFGUP1[8]  (.A(
        \ClockManagement_0/long_timer_0/count[9]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[8]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_4 ), .Y(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_6 ));
    XO1 \DUMP_0/dump_coder_0/para2_RNI4BP01[6]  (.A(
        \DUMP_0/count_0[6] ), .B(\DUMP_0/dump_coder_0/para2[6]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_3_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_1[0] ));
    IOPAD_BI \xd_pad[3]/U0/U0  (.D(\xd_pad[3]/U0/NET1 ), .E(
        \xd_pad[3]/U0/NET2 ), .Y(\xd_pad[3]/U0/NET3 ), .PAD(xd[3]));
    MX2 \top_code_0/relay_on_RNO_0[6]  (.A(\relay_on_c[6] ), .B(
        \GPMI_0_dataout[6] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_815 ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_0  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_14_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_20_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_5_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_0_Y ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]  (.D(
        \top_code_0_n_acqnum_2[9] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIQQUJ2[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_5[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_4[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_11[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_13[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[15]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[16]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_496 ));
    DFN1E1 \plusestate_0/PLUSETIME[2]  (.D(\top_code_0_plusedata[2] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[2]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[12]  (.D(
        \top_code_0_pd_pluse_data[12] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[12]_net_1 ));
    AX1C \DUMP_0/dump_timer_0/count_RNO_0[10]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_timer_0/count_c8 ), .C(\DUMP_0/count[10] ), .Y(
        \DUMP_0/dump_timer_0/count_n10_tz ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[4]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[4] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_4_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[4] ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_2  (.A(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .B(
        \timer_top_0/dataout[10] ), .C(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_2_Y ));
    IOIN_IB \xa_pad[9]/U0/U1  (.YIN(\xa_pad[9]/U0/NET1 ), .Y(\xa_c[9] )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_105  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_123_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_74_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_105_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[12]_net_1 ));
    NOR2B \DUMP_0/dump_state_0/cs4_0_o3  (.A(\DUMP_0/i_2[0] ), .B(
        state1ms_choice_0_reset_out), .Y(\DUMP_0/dump_state_0/cs4 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[19]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[20]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_508 ));
    IOPAD_IN \xa_pad[5]/U0/U0  (.PAD(xa[5]), .Y(\xa_pad[5]/U0/NET1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[4]  (.D(
        \DUMP_0/dump_coder_0/para2_4[4]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[4]_net_1 ));
    DFN1E1 \top_code_0/s_addchoice_0[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_0[0] ));
    AX1C \timer_top_0/timer_0/un2_timedata_I_35  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .C(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .Y(
        \timer_top_0/timer_0/I_35_1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[10]  (.A(
        \s_acq_change_0/s_stripnum_5[10] ), .B(
        \s_acq_change_0_s_stripnum[10] ), .S(\top_code_0_change[1] ), 
        .Y(\s_acq_change_0/N_66 ));
    NOR2A \scanstate_0/timecount_1_RNO[12]  (.A(\scanstate_0/N_70 ), 
        .B(\scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[12] ));
    DFN1E1 \scanstate_0/dectime[8]  (.D(\top_code_0_scandata[8] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[8]_net_1 ));
    MX2 \noisestate_0/soft_d_RNO_0  (.A(noisestate_0_soft_d), .B(
        \noisestate_0/CS[1]_net_1 ), .S(\noisestate_0/N_248 ), .Y(
        \noisestate_0/N_109 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[4]  (.D(
        \top_code_0_bri_datain[8] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[4] ));
    DFN1E1 \top_code_0/s_acqnum[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[10] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[8]_net_1 ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_3  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_2_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_1_Y ), .C(
        \timer_top_0/dataout[0] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_3_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_126  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_126_Y ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[5]  (.A(
        \s_acq_change_0/s_acqnum_5[5] ), .B(
        \s_acq_change_0_s_acqnum[5] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_75 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_7_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_7_net ));
    NOR2B \scanstate_0/rt_sw_RNO  (.A(\scanstate_0/N_111 ), .B(net_33), 
        .Y(\scanstate_0/rt_sw_RNO_2 ));
    DFN1 \scalestate_0/CS[20]  (.D(\scalestate_0/CS_RNO[20]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[20]_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[15]  (.D(
        \top_code_0_dds_configdata[14] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[15]_net_1 ));
    MX2 \bri_dump_sw_0/off_test_RNO_0  (.A(plusestate_0_off_test), .B(
        scalestate_0_off_test), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/off_test_5 ));
    IOTRI_OB_EB \k2_pad/U0/U1  (.D(k2_c), .E(VCC), .DOUT(
        \k2_pad/U0/NET1 ), .EOUT(\k2_pad/U0/NET2 ));
    DFN1 \top_code_0/relay_close[5]  (.D(
        \top_code_0/relay_close_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[5] ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[1]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[1] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[1]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m58  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_59 ));
    DFN1E1 \top_code_0/n_acqnum[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[2] ));
    OR2 \scalestate_0/CS_RNISQVB[21]  (.A(\scalestate_0/CS[1]_net_1 ), 
        .B(\scalestate_0/CS[21]_net_1 ), .Y(\scalestate_0/N_1201 ));
    XO1 \PLUSE_0/qq_coder_1/un1_qq_para2_NE_1[0]  (.A(
        \PLUSE_0/count_7[3] ), .B(\PLUSE_0/qq_para2[3] ), .C(
        \PLUSE_0/qq_coder_1/un1_qq_para2_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_1[0]_net_1 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[11]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[11] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_1[11] ));
    AO1B \scalestate_0/off_test_RNO_1  (.A(\scalestate_0/N_1262 ), .B(
        \scalestate_0/N_1263 ), .C(timer_top_0_clk_en_scale_0), .Y(
        \scalestate_0/N_1175 ));
    DFN1E1 \top_code_0/pd_pluse_data[8]  (.D(\GPMI_0_dataout[8] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[8] ));
    IOBI_IB_OB_EB \xd_pad[15]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[15] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[15]/U0/NET3 ), .DOUT(
        \xd_pad[15]/U0/NET1 ), .EOUT(\xd_pad[15]/U0/NET2 ), .Y(
        \xd_in[15] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[14]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c12 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n14 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_41_i ));
    DFN1E1 \top_code_0/state_1ms_data[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[0] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[13]_net_1 ));
    NOR2B \scalestate_0/dump_sustain_ctrl_RNO  (.A(
        \scalestate_0/N_744 ), .B(top_code_0_scale_rst_5), .Y(
        \scalestate_0/dump_sustain_ctrl_RNO_net_1 ));
    NOR2B \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_RNO  (.A(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_net_1 ), .B(net_27), .Y(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_RNO_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_2[4]  (.A(
        \state_1ms_0/M_DUMPTIME[4]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[4] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[4] ));
    DFN1E1 \plusestate_0/PLUSETIME[10]  (.D(\top_code_0_plusedata[10] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[10]_net_1 ));
    XO1 \DUMP_0/dump_coder_0/para3_RNIITV21[9]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_coder_0/para3[9]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_5[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[10]  (.A(
        \plusestate_0_timecount[10] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_254 ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[4]_net_1 ));
    OR3 \PLUSE_0/bri_coder_0/un2lto7_3  (.A(\PLUSE_0/count_2[5] ), .B(
        \PLUSE_0/count_2[7] ), .C(
        \PLUSE_0/bri_coder_0/un2lto7_1_net_1 ), .Y(
        \PLUSE_0/bri_coder_0/un2lto7_3_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_1  (.A(\ADC_c[9] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[8]_net_1 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[6]  (.D(
        \top_code_0_state_1ms_data[6] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[6]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIC4SG[11]  (.A(
        \DUMP_0/dump_coder_0/para3[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_11[0] ));
    NOR2A \scalestate_0/CS_RNIN85E[15]  (.A(\scalestate_0/N_1263 ), .B(
        \scalestate_0/CS[15]_net_1 ), .Y(\scalestate_0/N_1269 ));
    XOR2 \CAL_0/cal_div_0/count_RNIU6VJ[3]  (.A(
        \CAL_0/cal_div_0/count[3]_net_1 ), .B(\CAL_0/cal_para_out[3] ), 
        .Y(\CAL_0/cal_div_0/clear_n4_3 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_37_i ));
    NOR3C \scalestate_0/necount_LE_M_RNIPTOI  (.A(scalestate_0_ne_le), 
        .B(\scalestate_0/CS[12]_net_1 ), .C(
        \scalestate_0/necount_LE_M_net_1 ), .Y(
        \scalestate_0/timecount_12_sqmuxa_0 ));
    OR3A \top_code_0/pn_change_3_i_o2  (.A(\xa_c[6] ), .B(
        \top_code_0/N_137 ), .C(\top_code_0/N_140 ), .Y(
        \top_code_0/N_148 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[3]  (.D(\top_code_0_scaledatain[3] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[3]_net_1 ));
    NOR2B \bri_dump_sw_0/tetw_pluse_RNO  (.A(
        \bri_dump_sw_0/tetw_pluse_5 ), .B(net_27), .Y(
        \bri_dump_sw_0/tetw_pluse_RNO_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]  (.D(
        \top_code_0_n_acqnum_2[6] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]_net_1 ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[5]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_32 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[5] ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_3  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_4_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_1_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_8_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_3_Y ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m44_6 ));
    NOR2B \scalestate_0/timecount_ret_35_RNO_5  (.A(
        \scalestate_0/OPENTIME_TEL[9]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[9] ));
    CLKINT \GPMI_0/rst_n_module_0/rst_nr2_RNISUE8  (.A(
        \GPMI_0/rst_n_module_0/rst_nr2_net_1 ), .Y(net_27));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[7]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c6 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n7 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m41 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[18] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/SAND2_28_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net ), 
        .C(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_33_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_21_net ));
    NOR2B \scanstate_0/calctrl_RNO  (.A(\scanstate_0/N_131 ), .B(
        net_33), .Y(\scanstate_0/calctrl_RNO_net_1 ));
    NOR2B \scalestate_0/CS_RNO[16]  (.A(\scalestate_0/N_1229 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[16]_net_1 ));
    DFN1 \DUMP_OFF_0/off_on_timer_0/count[1]  (.D(
        \DUMP_OFF_0/off_on_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/count_3[1] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_9_inst  (.A(
        \sd_acq_top_0/count_3[6] ), .B(\sd_acq_top_0/count_3[7] ), .C(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ));
    DFN1 \DUMP_0/off_on_timer_1/count[1]  (.D(
        \DUMP_0/off_on_timer_1/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[1] ));
    IOPAD_TRI \Acq_clk_pad/U0/U0  (.D(\Acq_clk_pad/U0/NET1 ), .E(
        \Acq_clk_pad/U0/NET2 ), .PAD(Acq_clk));
    DFN1E1 \scalestate_0/PLUSETIME180[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[12]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[9]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[9]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/sd_sacq_state_0/cs[9]_net_1 ));
    OR3B \top_code_0/nstatechoice_3_i_o2_0  (.A(\xa_c[4] ), .B(
        \xa_c[7] ), .C(\top_code_0/N_139 ), .Y(\top_code_0/N_151 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_26  
        (.A(\s_acq_change_0_s_stripnum[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[4] )
        , .C(\s_acq_change_0_s_stripnum[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_26 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_12  
        (.A(\s_acq_change_0_s_stripnum[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .C(\s_acq_change_0_s_stripnum[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_12_0 ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ));
    DFN1 \scalestate_0/tetw_pluse  (.D(\scalestate_0/tetw_pluse_RNO_1 )
        , .CLK(GLA_net_1), .Q(scalestate_0_tetw_pluse));
    DFN1 \PLUSE_0/qq_state_0/stateover  (.D(
        \PLUSE_0/qq_state_0/stateover_RNO_0 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_0_stateover ));
    IOPAD_IN \xa_pad[2]/U0/U0  (.PAD(xa[2]), .Y(\xa_pad[2]/U0/NET1 ));
    OA1 \sd_acq_top_0/sd_sacq_state_0/cs_RNO[10]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_233 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_232 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[10] ));
    DFN1 \timer_top_0/timer_0/timedata[1]  (.D(
        \timer_top_0/timer_0/timedata_4[1] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[1]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m95  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_94 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_95 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_96 ));
    NOR3C \top_code_0/halfdata_1_sqmuxa_0_a2  (.A(\top_code_0/N_331 ), 
        .B(\top_code_0/N_334 ), .C(\top_code_0/N_329 ), .Y(
        \top_code_0/halfdata_1_sqmuxa ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[1]_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_4[9]  (.A(
        \state_1ms_0/S_DUMPTIME[9]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[9] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[9] ));
    DFN1 \syn_md_module_1/syn_md_0/count[3]  (.D(
        \syn_md_module_1/syn_md_0/count_RNO[3]_net_1 ), .CLK(GLA_net_1)
        , .Q(\syn_md_module_1/syn_md_0/count[3]_net_1 ));
    AND3 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_6  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] )
        );
    MX2 \state_1ms_0/soft_dump_RNO_0  (.A(state_1ms_0_soft_dump), .B(
        \state_1ms_0/N_255 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_152 ));
    OR3 \scalestate_0/timecount_ret_75_RNIPOAF  (.A(
        \scalestate_0/timecount_20_iv_9_reto[5] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[5] ), .C(
        \scalestate_0/timecount_cnst_m_reto[5] ), .Y(
        \scalestate_0_timecount[5] ));
    OR3 \scalestate_0/timecount_ret_50_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[17] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[17] ), .C(
        \scalestate_0/timecount_20_0_iv_2[17] ), .Y(
        \scalestate_0/timecount_20_0_iv_4[17] ));
    DFN1 \state_1ms_0/timecount[4]  (.D(
        \state_1ms_0/timecount_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[4] ));
    NOR2A \scalestate_0/intertodsp_RNO_3  (.A(
        \scalestate_0/CS[10]_net_1 ), .B(
        \scalestate_0/fst_lst_pulse_net_1 ), .Y(
        \scalestate_0/intertodsp_1_sqmuxa ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_163  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_88_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_1_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_163_Y ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_7  (.A(
        \timer_top_0/dataout[13] ), .B(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_8_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_7_Y ));
    OA1A \scalestate_0/CS_RNO[18]  (.A(\scalestate_0/N_1213 ), .B(
        \scalestate_0/CS[18]_net_1 ), .C(top_code_0_scale_rst_1), .Y(
        \scalestate_0/CS_RNO[18]_net_1 ));
    DFN1 \DDS_0/dds_state_0/w_clk_reg  (.D(
        \DDS_0/dds_state_0/w_clk_reg_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/w_clk_reg_net_1 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNO_0[15]  (.A(
        \ClockManagement_0/long_timer_0/count[14]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count_c13 ), .Y(
        \ClockManagement_0/long_timer_0/count_31_0 ));
    NOR2B \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_RNO  (.A(net_27), .B(xwe_c), 
        .Y(\GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_RNO_net_1 ));
    OR3A \top_code_0/relay_close_1_sqmuxa_0_o2_2  (.A(GPMI_0_code_en), 
        .B(\xa_c[18] ), .C(\top_code_0/un1_xa_30_0_o2_0_net_1 ), .Y(
        \top_code_0/N_137 ));
    MX2 \state_1ms_0/bri_cycle_RNO_0  (.A(state_1ms_0_bri_cycle), .B(
        \state_1ms_0/CS[5]_net_1 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_156 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_66  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_36_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_107_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_66_Y ));
    DFN1 \scalestate_0/necount[1]  (.D(
        \scalestate_0/necount_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[1]_net_1 ));
    DFN1 \nsctrl_choice_0/dumpon_ctr  (.D(
        \nsctrl_choice_0/dumpon_ctr_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_dumpon_ctr));
    OR3 \sd_acq_top_0/sd_sacq_state_0/en2_RNO_0  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_233 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_232 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_201 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/en2_0_0_o3_0 ));
    NOR3C \DUMP_0/off_on_timer_1/count_0_sqmuxa  (.A(
        \DUMP_0/dump_state_0_on_start ), .B(
        \DUMP_0/off_on_state_1_state_over ), .C(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ));
    DFN1E1 \top_code_0/noisedata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[5] ));
    AO1C \noisestate_0/CS_RNO_0[4]  (.A(\noisestate_0/CS[3]_net_1 ), 
        .B(timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[4] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[4]_net_1 ));
    NOR2B \nsctrl_choice_0/soft_d_RNO  (.A(\nsctrl_choice_0/soft_d_5 ), 
        .B(net_27), .Y(\nsctrl_choice_0/soft_d_RNO_0_net_1 ));
    AX1C \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_5_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[6] ));
    DFN1 \scanstate_0/CS[3]  (.D(\scanstate_0/CS_RNO_2[3] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[3]_net_1 ));
    DFN1 \ClockManagement_0/clk_10k_0/count[2]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[2] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[2]_net_1 ));
    NOR2 \top_code_0/s_addchoice_1_sqmuxa_0_a2_0  (.A(
        \top_code_0/N_144 ), .B(\top_code_0/N_164 ), .Y(
        \top_code_0/s_addchoice_1_sqmuxa_0_a2_0_net_1 ));
    INV \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBUBBLEA  (.A(
        n_acq_change_0_n_acq_start), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[1]  (.D(
        \DUMP_0/dump_coder_0/para4_4[1]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[1]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI4U1G[8]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[8]_net_1 ), 
        .B(\pd_pluse_top_0/count_0[8] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_8[0] ));
    DFN1E1 \scalestate_0/ACQ180_NUM[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[9]_net_1 ));
    NOR2B \DDS_0/dds_state_0/para_RNO_0[34]  (.A(
        \DDS_0/dds_state_0/para[35]_net_1 ), .B(
        \DDS_0/dds_state_0/N_534 ), .Y(\DDS_0/dds_state_0/N_524 ));
    PLLBA \ClockManagement_0/pllclk_0/Core  (.CLKA(OCX40MHz_c), .EXTFB(
        GND), .POWERDOWN(VCC), .GLA(GLA_net_1), .LOCK(), .GLB(
        \ClockManagement_0/pllclk_0_GLB ), .YB(), .GLC(), .YC(), 
        .OADIV0(GND), .OADIV1(GND), .OADIV2(GND), .OADIV3(GND), 
        .OADIV4(GND), .OAMUX0(GND), .OAMUX1(GND), .OAMUX2(VCC), 
        .DLYGLA0(GND), .DLYGLA1(GND), .DLYGLA2(GND), .DLYGLA3(GND), 
        .DLYGLA4(GND), .OBDIV0(VCC), .OBDIV1(VCC), .OBDIV2(GND), 
        .OBDIV3(GND), .OBDIV4(VCC), .OBMUX0(GND), .OBMUX1(VCC), 
        .OBMUX2(GND), .DLYYB0(GND), .DLYYB1(GND), .DLYYB2(GND), 
        .DLYYB3(GND), .DLYYB4(GND), .DLYGLB0(GND), .DLYGLB1(GND), 
        .DLYGLB2(GND), .DLYGLB3(GND), .DLYGLB4(GND), .OCDIV0(
        AFLSDF_GND), .OCDIV1(AFLSDF_GND), .OCDIV2(AFLSDF_GND), .OCDIV3(
        AFLSDF_GND), .OCDIV4(AFLSDF_GND), .OCMUX0(AFLSDF_GND), .OCMUX1(
        AFLSDF_GND), .OCMUX2(AFLSDF_GND), .DLYYC0(AFLSDF_GND), .DLYYC1(
        AFLSDF_GND), .DLYYC2(AFLSDF_GND), .DLYYC3(AFLSDF_GND), .DLYYC4(
        AFLSDF_GND), .DLYGLC0(AFLSDF_GND), .DLYGLC1(AFLSDF_GND), 
        .DLYGLC2(AFLSDF_GND), .DLYGLC3(AFLSDF_GND), .DLYGLC4(
        AFLSDF_GND), .FINDIV0(GND), .FINDIV1(VCC), .FINDIV2(GND), 
        .FINDIV3(GND), .FINDIV4(VCC), .FINDIV5(GND), .FINDIV6(GND), 
        .FBDIV0(GND), .FBDIV1(VCC), .FBDIV2(GND), .FBDIV3(GND), 
        .FBDIV4(VCC), .FBDIV5(GND), .FBDIV6(GND), .FBDLY0(GND), 
        .FBDLY1(GND), .FBDLY2(GND), .FBDLY3(GND), .FBDLY4(GND), 
        .FBSEL0(VCC), .FBSEL1(GND), .XDLYSEL(GND), .VCOSEL0(GND), 
        .VCOSEL1(GND), .VCOSEL2(VCC));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_2  (.A(\ADC_c[8] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_2 ));
    AO1 \scalestate_0/timecount_ret_51_RNO  (.A(
        \scalestate_0/OPENTIME[18]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[18] ), .Y(
        \scalestate_0/timecount_20_0_iv_0[18] ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_6_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_8_net ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[8] ));
    DFN1 \DUMP_ON_0/off_on_state_0/state_over  (.D(
        \DUMP_ON_0/off_on_state_0/N_9 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/off_on_state_0_state_over ));
    DFN1E1 \scalestate_0/NE_NUM[5]  (.D(\top_code_0_scaledatain[5] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[5]_net_1 ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_8  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_1_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_28_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_22_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_8_Y ));
    DFN1 \scalestate_0/CS[12]  (.D(\scalestate_0/CS_RNO[12]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_14  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_110_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_25_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_14_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m267  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_266 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_267 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_268 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIKOD81[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_4[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_15[0] ));
    AO1B \scalestate_0/tetw_pluse_RNO  (.A(\scalestate_0/N_1187 ), .B(
        scalestate_0_tetw_pluse), .C(top_code_0_scale_rst_1), .Y(
        \scalestate_0/tetw_pluse_RNO_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[8]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[10]_net_1 ));
    DFN1E1 \top_code_0/scandata[15]  (.D(\GPMI_0_dataout[15] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[15] ));
    NOR2B \state_1ms_0/timecount_RNO[14]  (.A(\state_1ms_0/N_81 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[14]_net_1 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[11]_net_1 ));
    AO1C \ClockManagement_0/long_timer_0/timeup_RNIUBFJ1  (.A(
        sigtimeup_c), .B(\ClockManagement_0/long_timer_0/clk_5K_en_1 ), 
        .C(\ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/counte ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[15]  (.D(
        \top_code_0_pd_pluse_data[15] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[15]_net_1 ));
    NOR2B \state1ms_choice_0/reset_out_RNO  (.A(
        \state1ms_choice_0/reset_out_5 ), .B(net_27), .Y(
        \state1ms_choice_0/reset_out_RNO_0_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[14]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[14] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[14] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[5]  (.A(
        \scalestate_0_strippluse[5] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[5] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[8]  (.A(
        \DDS_0/dds_state_0/para[8]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_282 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[8] ));
    DFN1E1 \plusestate_0/DUMPTIME[2]  (.D(\top_code_0_plusedata[2] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[2]_net_1 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ));
    XA1A \syn_md_module_1/syn_md_0/count_RNO_0[1]  (.A(
        \syn_md_module_1/syn_md_0/count[0]_net_1 ), .B(
        \syn_md_module_1/syn_md_0/count[1]_net_1 ), .C(
        \syn_md_module_1/syn_md_0/N_52 ), .Y(
        \syn_md_module_1/syn_md_0/count_RNO_0[1]_net_1 ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNISQPR1[1]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_1[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_4[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_7[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_11[0] ));
    NOR3A \top_code_0/un1_state_1ms_rst_n117_43_i_a2_1  (.A(
        \top_code_0/un1_state_1ms_rst_n117_43_i_a2_1_1_net_1 ), .B(
        \xa_c[6] ), .C(\top_code_0/N_137 ), .Y(\top_code_0/N_326 ));
    NOR2B \state_1ms_0/timecount_RNO_6[7]  (.A(
        \state_1ms_0/PLUSETIME[7]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[7] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m66  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_51 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_66 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[0] ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_72_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_24 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ));
    DFN1 \scanstate_0/calctrl  (.D(\scanstate_0/calctrl_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(scanstate_0_calctrl));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[4] ));
    NOR3C \PLUSE_0/qq_coder_0/i_RNO[1]  (.A(
        \PLUSE_0/qq_coder_0/i_0_4[1] ), .B(
        \PLUSE_0/qq_coder_0/un1_qq_para2_i[0] ), .C(
        \PLUSE_0/qq_coder_0/i_reg10_NE[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/i_RNO_6[1] ));
    OR3 \bridge_div_0/count_RNIDV0F1[4]  (.A(
        \bridge_div_0/count[5]_net_1 ), .B(
        \bridge_div_0/count[4]_net_1 ), .C(
        \bridge_div_0/un1_count_3[0] ), .Y(
        \bridge_div_0/un1_count_NE_0[0] ));
    NOR3B \pd_pluse_top_0/pd_pluse_coder_0/i_RNO[3]  (.A(net_27), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_i[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[3] ));
    XO1 \scalestate_0/fst_lst_pulse_RNO_7  (.A(
        \scalestate_0/necount[3]_net_1 ), .B(
        \scalestate_0/NE_NUM[3]_net_1 ), .C(
        \scalestate_0/fst_lst_pulse8_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_2 ));
    IOPAD_BI \xd_pad[13]/U0/U0  (.D(\xd_pad[13]/U0/NET1 ), .E(
        \xd_pad[13]/U0/NET2 ), .Y(\xd_pad[13]/U0/NET3 ), .PAD(xd[13]));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[2]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_187 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_173 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[2]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[10]  (.D(
        \DUMP_0/dump_coder_0/para5_4[10] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[10]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i16_mux ));
    DFN1E1 \scalestate_0/NE_NUM[4]  (.D(\top_code_0_scaledatain[4] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[4]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI6I0P[15]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[15]_net_1 ), .B(
        \sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_15[0] ));
    DFN1E1 \scalestate_0/ACQ90_NUM[9]  (.D(\top_code_0_scaledatain[9] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[9]_net_1 ));
    IOTRI_OB_EB \pd_pulse_en_pad/U0/U1  (.D(pd_pulse_en_c), .E(VCC), 
        .DOUT(\pd_pulse_en_pad/U0/NET1 ), .EOUT(
        \pd_pulse_en_pad/U0/NET2 ));
    NOR2B \nsctrl_choice_0/rt_sw_RNO  (.A(\nsctrl_choice_0/rt_sw_5 ), 
        .B(net_27), .Y(\nsctrl_choice_0/rt_sw_RNO_0_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[3]  (.A(
        \scanstate_0_timecount[3] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_226 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIJA8G[3]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11 ), 
        .B(\s_acq_change_0_s_stripnum[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_3 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIG2DH[19]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[19]_net_1 ), .B(
        \sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_19[0] ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/count_RNO_0[3]  (.A(
        \DSTimer_0/dump_sustain_timer_0/count[2]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count_c1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_7_0 ));
    DFN1E1 \top_code_0/n_acqnum[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[8] ));
    IOBI_IB_OB_EB \xd_pad[9]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[9] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[9]/U0/NET3 ), .DOUT(\xd_pad[9]/U0/NET1 ), .EOUT(
        \xd_pad[9]/U0/NET2 ), .Y(\xd_in[9] ));
    DFN1 \DUMP_0/dump_coder_0/i[4]  (.D(
        \DUMP_0/dump_coder_0/i_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i[4] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[0]  (.D(
        \top_code_0_state_1ms_data[0] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[0]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[9]  (.A(
        \scanstate_0_timecount[9] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_201 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i2_mux ));
    DFN1E1 \top_code_0/pn_change  (.D(\top_code_0/N_92 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pn_change));
    DFN1E1 \top_code_0/scandata[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[9] ));
    DFN1E1 \state_1ms_0/PLUSETIME[14]  (.D(
        \top_code_0_state_1ms_data[14] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[14]_net_1 ));
    AO1C \state_1ms_0/CS_RNO_0[2]  (.A(\state_1ms_0/CS[1]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[2] ));
    OR3A \ClockManagement_0/clk_div500_0/count_RNO[0]  (.A(net_27), .B(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .C(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_partial_sum[0] )
        , .Y(\ClockManagement_0/clk_div500_0/count_5[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m41_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[18] ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_4  (.A(
        \scalestate_0/necount[2]_net_1 ), .B(
        \scalestate_0/NE_NUM[2]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_4_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[27]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[28]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_476 ));
    NOR3B \state_1ms_0/PLUSETIME_1_sqmuxa_0_a2  (.A(
        \top_code_0_state_1ms_lc[0] ), .B(\state_1ms_0/N_17 ), .C(
        \top_code_0_state_1ms_lc[1] ), .Y(
        \state_1ms_0/PLUSETIME_1_sqmuxa ));
    DFN1E1 \scalestate_0/timecount_ret_31  (.D(
        \scalestate_0/timecount_20_iv_3[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_3_reto[4] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[1]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n1 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[15]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_43 ), .Y(
        \timer_top_0/timer_0/timedata_4[15] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_121  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_121_Y ));
    DFN1E1 \scalestate_0/CUTTIME90[17]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[17]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[7]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c6 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[7] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n7 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[0]  (.A(
        \Signal_Noise_Acq_0/un1_signal_acq_0[0] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_0_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[0] ));
    XO1 \DUMP_0/dump_coder_0/para4_RNIO6551[2]  (.A(
        \DUMP_0/count_1[2] ), .B(\DUMP_0/dump_coder_0/para4[2]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_1_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_3[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m26  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_23 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_26 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_27 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[3]  (.A(
        \Signal_Noise_Acq_0/un1_signal_acq_0[3] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_3_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[3] ));
    MX2 \scalestate_0/necount_RNO_0[1]  (.A(\scalestate_0/necount1[1] )
        , .B(\scalestate_0/necount[1]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_731 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[8]  (.A(
        \top_code_0_s_acqnum_2[8] ), .B(\scalestate_0_s_acqnum[8] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[8] ));
    NOR3C \scalestate_0/timecount_ret_88_RNO_0  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[10]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[10] ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[11]  (.A(\scalestate_0/N_558 ), 
        .B(top_code_0_scale_rst_4), .Y(
        \scalestate_0/s_acqnum_1_RNO[11]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_53  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_53_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_68  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_149_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_138_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_68_Y ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[3]  (.D(
        \top_code_0_pd_pluse_data[3] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[3]_net_1 ));
    DFN1E1 \scalestate_0/ACQTIME[3]  (.D(\top_code_0_scaledatain_0[3] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[3]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[21]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[21]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[21] ));
    MX2 \state_1ms_0/dump_start_RNO_0  (.A(state_1ms_0_dump_start), .B(
        \state_1ms_0/N_256 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_87 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[1]  (.A(
        \scanstate_0_timecount[1] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_236 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_45  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[2] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[3] )
        );
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIO1QF[3]  (.A(
        \sd_acq_top_0/count_10[3] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[3]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_0[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_7[0] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m57  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[3]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_58_i ));
    NOR2B \scalestate_0/timecount_ret_69_RNO_1  (.A(
        \scalestate_0/OPENTIME[15]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[15] ));
    DFN1 \top_code_0/scale_rst_4  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_4));
    DFN1 \DUMP_ON_0/off_on_timer_0/count[4]  (.D(
        \DUMP_ON_0/off_on_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/count_5[4] ));
    AND3 \CAL_0/cal_div_0/un3_count_I_8  (.A(
        \CAL_0/cal_div_0/count[0]_net_1 ), .B(
        \CAL_0/cal_div_0/count[1]_net_1 ), .C(
        \CAL_0/cal_div_0/count[2]_net_1 ), .Y(\CAL_0/cal_div_0/N_4 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[9]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c8 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n9 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ));
    DFN1E1 \scalestate_0/ACQTIME[9]  (.D(\top_code_0_scaledatain[9] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[9]_net_1 ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[10]  (.A(
        \sd_acq_top_0/count_1[8] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[8]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_2[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_4[10] ));
    DFN1 \scanstate_0/CS[6]  (.D(\scanstate_0/CS_RNO_2[6] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[6]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_55  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[28] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[13] ), .C(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .Y(
        \timer_top_0/timer_0/N_4 ));
    DFN1E1 \top_code_0/n_s_ctrl_0  (.D(\top_code_0/N_76 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_n_s_ctrl_0));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i6_mux ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i20_mux ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[5]  (.D(
        \top_code_0_state_1ms_data[5] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[5]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_19  (.D(
        \scalestate_0/timecount_20_iv_3[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_3_reto[8] ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIKMS51[11]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3 ), .B(
        \s_acq_change_0_s_stripnum[11] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_11 ));
    DFN1E1 \top_code_0/cal_data[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[0] ));
    MX2 \plusestate_0/timecount_1_RNO_0[10]  (.A(
        \plusestate_0/DUMPTIME[10]_net_1 ), .B(
        \plusestate_0/PLUSETIME[10]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_81 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[11]  (.A(
        \noisestate_0_timecount[11] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_195 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_41_i ));
    NOR2A \scalestate_0/timecount_ret_71_RNO_4  (.A(
        \scalestate_0/CUTTIME90[15]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[15] ));
    AO1 \scalestate_0/timecount_ret_1_RNO_1  (.A(
        \scalestate_0/CUTTIME180[5]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[5] ), .Y(
        \scalestate_0/timecount_20_iv_2[5] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[21]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[21]_net_1 ));
    AO1D \scalestate_0/CS_0_RNIAQA34[11]  (.A(\scalestate_0/N_1153_1 ), 
        .B(\scalestate_0/CS_0[11]_net_1 ), .C(
        \scalestate_0/un1_CS6_26_0 ), .Y(\scalestate_0/un1_CS6_26 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[0]  (.D(
        \DUMP_0/dump_coder_0/para4_4[0]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[0]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m265  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_266 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[32]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[32]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_313 ));
    NOR3B \scalestate_0/DUMPTIME_1_sqmuxa_0_a2  (.A(
        \scalestate_0/N_61 ), .B(\scalestate_0/N_60 ), .C(
        \top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/DUMPTIME_1_sqmuxa ));
    MX2B \scanstate_0/timecount_1_RNO[9]  (.A(\scanstate_0/N_67 ), .B(
        \scanstate_0/N_196 ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[9] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[5]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[6]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_323 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_129  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_129_Y ));
    NOR2 \top_code_0/relay_on_1_sqmuxa_0_a2_0  (.A(\xa_c[0] ), .B(
        \xa_c[1] ), .Y(\top_code_0/N_329 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[7]  (.A(
        \scalestate_0_timecount[7] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_208 ));
    DFN1 \timer_top_0/state_switch_0/dataout[3]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[3]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[3] ));
    MX2 \scalestate_0/necount_RNO_0[6]  (.A(\scalestate_0/necount1[6] )
        , .B(\scalestate_0/necount[6]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_736 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[4]  (.A(
        \s_acq_change_0/s_stripnum_5[4] ), .B(
        \s_acq_change_0_s_stripnum[4] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_60 ));
    NOR2B \top_code_0/un1_xa_8_16_i_i_o3_i_a2  (.A(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_5_net_1 ), .B(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_4_net_1 ), .Y(
        \top_code_0/N_13 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[5]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[5] ));
    DFN1 \s_acq_change_0/s_acqnum[3]  (.D(
        \s_acq_change_0/s_acqnum_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[3] ));
    OR3 \scalestate_0/timecount_ret_28_RNO  (.A(
        \scalestate_0/S_DUMPTIME_m[1] ), .B(
        \scalestate_0/timecount_20_iv_1[1] ), .C(
        \scalestate_0/timecount_20_iv_7[1] ), .Y(
        \scalestate_0/timecount_20_iv_9[1] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_8_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_8_net ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[20]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[20]_net_1 ));
    NOR3B \DUMP_ON_0/off_on_coder_0/i_RNO_0[1]  (.A(
        \DUMP_ON_0/count_5[4] ), .B(\DUMP_ON_0/count_5[2] ), .C(
        \DUMP_ON_0/count_5[3] ), .Y(
        \DUMP_ON_0/off_on_coder_0/i_0_2[1] ));
    XOR2 \scalestate_0/necount_inc_0/FOR2_8_inst  (.A(
        \scalestate_0/necount_inc_0/Rcout_10_net ), .B(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/necount1[10] ));
    AO1A \noisestate_0/dumpon_ctr_RNO_0  (.A(
        \noisestate_0/CS[2]_net_1 ), .B(noisestate_0_dumpon_ctr), .C(
        \noisestate_0/CS[1]_net_1 ), .Y(\noisestate_0/N_130 ));
    IOPAD_IN \ADC_pad[0]/U0/U0  (.PAD(ADC[0]), .Y(\ADC_pad[0]/U0/NET1 )
        );
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIQ58R[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_6[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_7[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_11[0] ));
    NOR2B \CAL_0/cal_div_0/count_RNIMK654[1]  (.A(
        \CAL_0/cal_div_0/clear_n ), .B(scanstate_0_calctrl), .Y(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m110  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_109 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_110 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_111 ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_48_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[5] )
        );
    DFN1 \DUMP_0/off_on_timer_0/count[1]  (.D(
        \DUMP_0/off_on_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_2[1] ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[1] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_70_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n5 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5]/Y ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_19  (.A(
        \top_code_0_sigtimedata[2] ), .B(
        \ClockManagement_0/long_timer_0/count[2]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_2 ));
    AND3 \CAL_0/cal_div_0/un3_count_I_13  (.A(
        \CAL_0/cal_div_0/DWACT_FINC_E[0] ), .B(
        \CAL_0/cal_div_0/count[3]_net_1 ), .C(
        \CAL_0/cal_div_0/count[4]_net_1 ), .Y(\CAL_0/cal_div_0/N_2 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[16]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[16]_net_1 ));
    AO1 \scalestate_0/necount_cmp_1/AO1_0  (.A(
        \scalestate_0/necount_cmp_1/AND2_0_Y ), .B(
        \scalestate_0/necount_cmp_1/NAND3A_1_Y ), .C(
        \scalestate_0/necount_cmp_1/NOR3_0_Y ), .Y(
        \scalestate_0/necount_cmp_1/AO1_0_Y ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_4  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_19_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_23_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_2_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_4_Y ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[11]  (.D(
        \DUMP_0/dump_coder_0/para2_4[11]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[11]_net_1 ));
    MX2 \scalestate_0/necount_RNO_0[8]  (.A(\scalestate_0/necount1[8] )
        , .B(\scalestate_0/necount[8]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_738 ));
    OR2 \pd_pluse_top_0/pd_pluse_state_0/cs_RNIOV4D[3]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[3]_net_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_166 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m222  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_221 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_222 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_223 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[12]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNINUII[7]  (.A(
        \DUMP_0/dump_coder_0/para4[7]_net_1 ), .B(\DUMP_0/count_0[7] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_7[0] ));
    AO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_35  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[1] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[0] )
        );
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m72  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_73 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_23  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_23_Y ));
    AND2A \PLUSE_0/bri_coder_0/half_0_I_12  (.A(\PLUSE_0/count_2[7] ), 
        .B(\PLUSE_0/half_para[7] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[5] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i14_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[6]_net_1 ));
    IOPAD_TRI \ddsfqud_pad/U0/U0  (.D(\ddsfqud_pad/U0/NET1 ), .E(
        \ddsfqud_pad/U0/NET2 ), .PAD(ddsfqud));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_85  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_85_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_89  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_40_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_92_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_89_Y ));
    NOR2B \scalestate_0/timecount_ret_2_RNO_4  (.A(
        \scalestate_0/CUTTIME180[6]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[6] ));
    DFN1E1 \scalestate_0/ACQTIME[15]  (.D(\top_code_0_scaledatain[15] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[15]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[3]  (.D(\top_code_0_scaledatain[3] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[3]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m45_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] ));
    IOBI_IB_OB_EB \xd_pad[3]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[3] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[3]/U0/NET3 ), .DOUT(\xd_pad[3]/U0/NET1 ), .EOUT(
        \xd_pad[3]/U0/NET2 ), .Y(\xd_in[3] ));
    DFN1E1 \scalestate_0/M_NUM[6]  (.D(\top_code_0_scaledatain[6] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[6]_net_1 ));
    IOPAD_TRI \relay_close_pad[6]/U0/U0  (.D(
        \relay_close_pad[6]/U0/NET1 ), .E(\relay_close_pad[6]/U0/NET2 )
        , .PAD(relay_close[6]));
    DFN1 \DDS_0/dds_state_0/cs[7]  (.D(\DDS_0/dds_state_0/N_80 ), .CLK(
        GLA_net_1), .Q(\DDS_0/dds_state_0/cs[7]_net_1 ));
    NOR2B \scalestate_0/necount_LE_M_RNO  (.A(
        \scalestate_0/necount_LE_M_1 ), .B(top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_LE_M_RNO_net_1 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c2 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n4 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNICN6B[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[8]_net_1 ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_8[0] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_9_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_9_net ));
    DFN1E0 \DDS_0/dds_state_0/para[1]  (.D(\DDS_0/dds_state_0/N_46 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[1]_net_1 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[15]  (.D(
        \ClockManagement_0/long_timer_0/count_n15 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[15]_net_1 ));
    AO1 \PLUSE_0/bri_state_0/cs_RNO_1[3]  (.A(
        \PLUSE_0/bri_state_0/N_144 ), .B(clk_4f_en), .C(
        \PLUSE_0/bri_state_0/csse_2_0_0 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_1 ));
    IOIN_IB \xa_pad[5]/U0/U1  (.YIN(\xa_pad[5]/U0/NET1 ), .Y(\xa_c[5] )
        );
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m191  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_192 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m41_4 ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/data[2]  (.D(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[2]_net_1 ), .CLK(
        GLA_net_1), .Q(\DSTimer_0/dump_sustain_timer_0/data[2]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_38_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m44_2 ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_i_a2_0  (
        .A(\top_code_0_sd_sacq_choice[3] ), .B(
        \top_code_0_sd_sacq_choice[1] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_i_a2_0_net_1 )
        );
    XOR2 \CAL_0/cal_div_0/un3_count_I_5  (.A(
        \CAL_0/cal_div_0/count[0]_net_1 ), .B(
        \CAL_0/cal_div_0/count[1]_net_1 ), .Y(\CAL_0/cal_div_0/I_5 ));
    MX2 \top_code_0/relay_on_RNO_0[9]  (.A(\relay_on_c[9] ), .B(
        \GPMI_0_dataout[9] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_818 ));
    DFN1 \timer_top_0/state_switch_0/dataout[17]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[17]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[17] ));
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_41 ), .B(
        n_acq_change_0_n_rst_n), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_net_1 ));
    NOR2A \scalestate_0/timecount_ret_47_RNO_3  (.A(
        \scalestate_0/CUTTIME90[16]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[16] ));
    XOR2 \CAL_0/cal_div_0/un3_count_I_9  (.A(\CAL_0/cal_div_0/N_4 ), 
        .B(\CAL_0/cal_div_0/count[3]_net_1 ), .Y(\CAL_0/cal_div_0/I_9 )
        );
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m1  (.A(
        \top_code_0_n_divnum_0[5] ), .B(\top_code_0_n_divnum_0[0] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_i ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/data[3]  (.D(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[3]_net_1 ), .CLK(
        GLA_net_1), .Q(\DSTimer_0/dump_sustain_timer_0/data[3]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[1] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_68_i ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m47_6 ));
    XO1 \CAL_0/cal_div_0/count_RNIQBU71[2]  (.A(
        \CAL_0/cal_para_out[2] ), .B(\CAL_0/cal_div_0/count[2]_net_1 ), 
        .C(\CAL_0/cal_div_0/clear_n4_3 ), .Y(
        \CAL_0/cal_div_0/clear_n4_NE_1 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_5  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_5_1 ));
    AO1C \plusestate_0/timecount_1_RNO_1[1]  (.A(
        \plusestate_0/CS[3]_net_1 ), .B(\plusestate_0/CS_i[0]_net_1 ), 
        .C(top_code_0_pluse_rst_0), .Y(\plusestate_0/N_245 ));
    DFN1E1 \scalestate_0/timecount_ret_20  (.D(
        \scalestate_0/timecount_20_iv_8[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[8] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[11]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[11] ));
    DFN1 \scalestate_0/s_acqnum_1[5]  (.D(
        \scalestate_0/s_acqnum_1_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[5] ));
    DFN1E1 \noisestate_0/timecount_1[0]  (.D(
        \noisestate_0/timecount_5[0] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[0] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[10]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[10] ));
    NOR3B \top_code_0/change_1_sqmuxa_0_a2  (.A(\top_code_0/N_331 ), 
        .B(\top_code_0/N_329 ), .C(\top_code_0/N_154 ), .Y(
        \top_code_0/change_1_sqmuxa ));
    DFN1 \ClockManagement_0/clk_div500_0/clk_5K  (.D(
        \ClockManagement_0/clk_div500_0/clk_5K_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(\ClockManagement_0/clk_div500_0_clk_5K ));
    DFN1E1 \top_code_0/s_addchoice[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice[2] ));
    NOR3A \top_code_0/k1_RNO_4  (.A(\xa_c[7] ), .B(\xa_c[18] ), .C(
        \xa_c[1] ), .Y(\top_code_0/un1_state_1ms_rst_n117_5_i_a2_2 ));
    NOR3A \syn_md_module_1/syn_md_0/syn_md_out_RNO  (.A(
        top_code_0_scale_rst_0), .B(\syn_md_module_1/syn_md_0/N_30 ), 
        .C(\syn_md_module_1/syn_md_0/N_31 ), .Y(
        \syn_md_module_1/syn_md_0/N_14 ));
    DFN1E1 \top_code_0/bri_datain[15]  (.D(\GPMI_0_dataout[15] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[15] ));
    DFN1 \scalestate_0/strippluse[0]  (.D(
        \scalestate_0/strippluse_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[0] ));
    NOR3A \scalestate_0/necount_cmp_1/NOR3A_2  (.A(
        \scalestate_0/necount_cmp_1/OR2A_1_Y ), .B(
        \scalestate_0/necount_cmp_1/AO1C_0_Y ), .C(
        \scalestate_0/NE_NUM[0]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/NOR3A_2_Y ));
    NOR2A \PLUSE_0/bri_state_0/cs_RNO_3[3]  (.A(\PLUSE_0/i_1[4] ), .B(
        \PLUSE_0/i_3[3] ), .Y(\PLUSE_0/bri_state_0/csse_2_0_a4_2_5 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[12]  (.D(
        \top_code_0_state_1ms_data[12] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[12]_net_1 ));
    NOR2B \pd_pluse_top_0/pd_pluse_state_0/un1_state_initial_0_o5  (.A(
        \pd_pluse_top_0/i_6[0] ), .B(net_27), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ));
    MX2 \scanstate_0/timecount_1_RNO[7]  (.A(\scanstate_0/N_65 ), .B(
        \scanstate_0/timecount_cnst[4] ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[7] ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_4[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_3[10] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_14[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_18[10] ));
    DFN1E1 \top_code_0/sd_sacq_data[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[13] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_24  (.A(
        \timer_top_0/dataout[12] ), .B(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_24_Y ));
    DFN1E1 \top_code_0/nstateload  (.D(\top_code_0/N_80 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_nstateload));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_46  (.A(
        \timer_top_0/timer_0/N_7 ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .Y(
        \timer_top_0/timer_0/I_46 ));
    DFN1 \timer_top_0/state_switch_0/dataout[15]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[15]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[15] ));
    DFN1E1 \top_code_0/s_addchoice_1[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_1[1] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m302  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] ), .C(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_303 ));
    MX2 \scalestate_0/strippluse_RNO_0[5]  (.A(
        \scalestate_0/strippluse_6[5] ), .B(
        \scalestate_0_strippluse[5] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_564 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_37  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_50_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[2] )
        );
    NOR2 \plusestate_0/CS_RNIHRHP[3]  (.A(\plusestate_0/CS[3]_net_1 ), 
        .B(\plusestate_0/CS[4]_net_1 ), .Y(\plusestate_0/N_301 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_41  (.A(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[14]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[9] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ));
    DFN1E1 \scalestate_0/OPENTIME[19]  (.D(\top_code_0_scaledatain[3] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1681 ), .Q(
        \scalestate_0/OPENTIME[19]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_6[11]  (.A(
        \state_1ms_0/PLUSETIME[11]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[11] ));
    DFN1 \PLUSE_0/qq_state_0/cs[2]  (.D(
        \PLUSE_0/qq_state_0/cs_RNO_1[2]_net_1 ), .CLK(GLA_net_1), .Q(
        Q3Q6_c));
    AO1A \scalestate_0/timecount_20_iv_4[11]  (.A(
        \scalestate_0/N_1069 ), .B(\scalestate_0/CUTTIME90[11]_net_1 ), 
        .C(\scalestate_0/CUTTIMEI90_m[11] ), .Y(
        \scalestate_0/timecount_20_iv_4[11]_net_1 ));
    OA1A \scalestate_0/necount_cmp_1/OA1A_0  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/NE_NUM[9]_net_1 ), .C(
        \scalestate_0/NE_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OA1A_0_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[14]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[15]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_464 ));
    MX2 \scalestate_0/rt_sw_RNO_0  (.A(scalestate_0_rt_sw), .B(
        \scalestate_0/un1_CS_34 ), .S(\scalestate_0/N_1259 ), .Y(
        \scalestate_0/N_544 ));
    NOR3A \top_code_0/n_rd_en_RNO_1  (.A(\top_code_0/N_329 ), .B(
        \top_code_0/N_154 ), .C(\top_code_0/N_152 ), .Y(
        \top_code_0/N_282 ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[1]_net_1 ));
    DFN1 \PLUSE_0/qq_state_1/stateover  (.D(
        \PLUSE_0/qq_state_1/stateover_RNO_1 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_1_stateover ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[7]  (.A(
        \PLUSE_0/bri_state_0/cs_i_0[7] ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[6] ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_0[7] ));
    NOR2B \state_1ms_0/timecount_RNO[5]  (.A(\state_1ms_0/N_72 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[5]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[2]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[2] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[2]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[1]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[2]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_281 ));
    XA1C \ClockManagement_0/long_timer_0/timeup_RNO_11  (.A(
        \ClockManagement_0/long_timer_0/count[11]_net_1 ), .B(
        \top_code_0_sigtimedata[11] ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_13 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_1 ));
    NOR3B \scalestate_0/OPENTIME_TEL_560_e  (.A(\scalestate_0/N_64 ), 
        .B(\scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0_0[0] ), 
        .Y(\scalestate_0/N_1773 ));
    DFN1E1 \noisestate_0/dectime[4]  (.D(\top_code_0_noisedata[4] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[4]_net_1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[5]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c4 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n5 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m237  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_236 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_237 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_238 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI5L7O[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c2 ));
    NOR3C \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_2_i ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[7]  (.A(
        \top_code_0_dumpdata_0[7] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[7]_net_1 ));
    DFN1E1 \state_1ms_0/PLUSETIME[13]  (.D(
        \top_code_0_state_1ms_data[13] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[13]_net_1 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[3]  (.D(
        \top_code_0_state_1ms_data[3] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[3]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[5]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[5] ));
    XO1 \PLUSE_0/qq_coder_1/un1_qq_para2_NE_2[0]  (.A(
        \PLUSE_0/count_7[1] ), .B(\PLUSE_0/qq_para2[1] ), .C(
        \PLUSE_0/qq_coder_1/un1_qq_para2_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_2[0]_net_1 ));
    OR2A \scalestate_0/necount_cmp_0/OR2A_1  (.A(
        \scalestate_0/M_NUM[2]_net_1 ), .B(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_1_Y ));
    DFN1E1 \noisestate_0/timecount_1[4]  (.D(
        \noisestate_0/timecount_5[4] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[4] ));
    NOR2A \DDS_0/dds_state_0/cs_RNO[8]  (.A(\DDS_0/dds_state_0/N_223 ), 
        .B(\DDS_0/dds_state_0/N_451 ), .Y(
        \DDS_0/dds_state_0/cs_RNO[8]_net_1 ));
    IOIN_IB \xa_pad[2]/U0/U1  (.YIN(\xa_pad[2]/U0/NET1 ), .Y(\xa_c[2] )
        );
    NOR2B \s_acq_change_0/s_stripnum_RNO[1]  (.A(\s_acq_change_0/N_57 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[1]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m63  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_62 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_63 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_64 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[4]_net_1 ));
    NOR2B \top_code_0/plusedata_1_sqmuxa_0_a2_0  (.A(
        \top_code_0/N_332 ), .B(\top_code_0/N_333 ), .Y(
        \top_code_0/N_340 ));
    AO1C \state_1ms_0/CS_RNO_0[6]  (.A(\state_1ms_0/CS[5]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[6] ));
    OR2B \scalestate_0/CS_RNIBR8M[16]  (.A(\scalestate_0/CS[16]_net_1 )
        , .B(\scalestate_0/N_1196 ), .Y(\scalestate_0/N_1181 ));
    AO1C \noisestate_0/CS_RNO_0[2]  (.A(\noisestate_0/CS[1]_net_1 ), 
        .B(timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[2] ));
    OR3 \DUMP_0/dump_coder_0/para5_RNIC7AK2[0]  (.A(
        \DUMP_0/dump_coder_0/un1_count_10[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_0[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_8[0] ));
    DFN1E1 \top_code_0/halfdata[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[1] ));
    NOR2B \scalestate_0/timecount_ret_66_RNO_1  (.A(
        \scalestate_0/OPENTIME[14]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[14] ));
    OR3 \scalestate_0/timecount_ret_26_RNIRFA1  (.A(
        \scalestate_0/timecount_20_iv_9_reto[11] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[11] ), .C(
        \scalestate_0/timecount_11_sqmuxa_m_reto ), .Y(
        \scalestate_0_timecount[11] ));
    NOR3B \top_code_0/relay_on_1_sqmuxa_0_a2_0_0  (.A(
        \top_code_0/N_337 ), .B(\top_code_0/N_329 ), .C(
        \top_code_0/N_154 ), .Y(
        \top_code_0/relay_on_1_sqmuxa_0_a2_0_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[9]  (.A(
        \state_1ms_0/PLUSECYCLE[9]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[9] ));
    MX2 \scanstate_0/timecount_1_RNO_0[14]  (.A(
        \scanstate_0/acqtime[14]_net_1 ), .B(
        \scanstate_0/dectime[14]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_72 ));
    DFN1 \PLUSE_0/qq_timer_1/count[1]  (.D(
        \PLUSE_0/qq_timer_1/count_n1 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_7[1] ));
    NOR3 \topctrlchange_0/sw_acq2_RNO_2  (.A(\top_code_0_change_0[0] ), 
        .B(\top_code_0_change[1] ), .C(nsctrl_choice_0_sw_acq2), .Y(
        \topctrlchange_0/sw_acq2in1_i_m ));
    IOPAD_IN \xa_pad[15]/U0/U0  (.PAD(xa[15]), .Y(\xa_pad[15]/U0/NET1 )
        );
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNIENBF1[4]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c2 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c4 ));
    AO1C \noisestate_0/CS_RNO_0[5]  (.A(\noisestate_0/CS[4]_net_1 ), 
        .B(timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[5] ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_9  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_7_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_4_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_26_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_9_Y ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[9]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[9] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[14]_net_1 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[10]  (.D(
        \ClockManagement_0/long_timer_0/count_n10 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[10]_net_1 ));
    DFN1E1 \top_code_0/plusedata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[6] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[18]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[18]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_502 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_14  (.A(
        \timer_top_0/timer_0/N_18 ), .B(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .Y(
        \timer_top_0/timer_0/I_14_1 ));
    NOR2B \scalestate_0/CS_RNO[12]  (.A(\scalestate_0/N_1226 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[12]_net_1 ));
    DFN1E1 \scalestate_0/ACQTIME[6]  (.D(\top_code_0_scaledatain[6] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[6]_net_1 ));
    NOR2B \noisestate_0/CS_i_0_RNIIEDN[0]  (.A(\noisestate_0/CS_li[0] )
        , .B(\noisestate_0/N_250 ), .Y(\noisestate_0/N_248 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[5]_net_1 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[20]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_59 ), .Y(
        \timer_top_0/timer_0/timedata_4[20] ));
    NOR2B \plusestate_0/off_test_RNO  (.A(\plusestate_0/N_141 ), .B(
        top_code_0_pluse_rst), .Y(\plusestate_0/off_test_RNO_0_net_1 ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[7]  (.A(
        \DUMP_0/dump_timer_0/count_c6 ), .B(\DUMP_0/count_0[7] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n7 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m42_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[17] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI3I6T[13]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[13]_net_1 ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_13[0] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_5  (.A(\xd_in[9] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[9] ));
    AO1C \scanstate_0/CS_RNO_0[3]  (.A(\scanstate_0/CS[2]_net_1 ), .B(
        timer_top_0_clk_en_scan), .C(net_33_0), .Y(
        \scanstate_0/CS_srsts_i_0[3] ));
    DFN1E1 \scalestate_0/M_NUM[9]  (.D(\top_code_0_scaledatain[9] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[9]_net_1 ));
    DFN1E1 \plusestate_0/timecount_1[3]  (.D(
        \plusestate_0/timecount_5[3] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[3] ));
    MX2A \scalestate_0/sw_acq1_RNO_0  (.A(\scalestate_0/un1_CS_20 ), 
        .B(scalestate_0_sw_acq1), .S(\scalestate_0/un1_CS6_34 ), .Y(
        \scalestate_0/N_542 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m199  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_198 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_199 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_200 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/dataout[14]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[14] ), .B(
        top_code_0_n_s_ctrl_1), .Y(\Signal_Noise_Acq_0_dataout[14] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_6  (.A(\xd_in[8] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[8] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[10]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[9] ), 
        .Y(\DDS_0/dds_state_0/N_290 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[10]  (.A(
        \top_code_0_dumpdata_0[10] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[10]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[5]  (.D(\GPMI_0_dataout[5] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[5] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m47_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] ));
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_4  (.A(
        \scalestate_0/necount_cmp_1/NOR3A_2_Y ), .B(
        \scalestate_0/necount_cmp_1/OR2A_4_Y ), .C(
        \scalestate_0/necount_cmp_1/NAND3A_5_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_4_Y ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[1]  (.A(
        \scalestate_0/s_acqnum_7[1] ), .B(\scalestate_0_s_acqnum[1] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_548 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[11]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i6_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_160  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_160_Y ));
    OR2 \PLUSE_0/qq_coder_1/i_reg10_NE[0]  (.A(
        \PLUSE_0/qq_coder_1/i_reg10_NE_3[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_1/i_reg10_NE_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_NE[0]_net_1 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[15]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[15] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count[15] ));
    DFN1 \timer_top_0/timer_0/timedata[19]  (.D(
        \timer_top_0/timer_0/timedata_4[19] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[19]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m23  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_24 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_114  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_114_Y ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[8]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c6 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n8 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[3]  (.D(
        \top_code_0_pd_pluse_data[3] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m218  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_215 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_218 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_219 ));
    DFN1 \nsctrl_choice_0/rt_sw  (.D(
        \nsctrl_choice_0/rt_sw_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_rt_sw));
    DFN1E1 \scalestate_0/M_NUM[3]  (.D(\top_code_0_scaledatain_0[3] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[3]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[8]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[11]  (.A(
        \noisestate_0/acqtime[11]_net_1 ), .B(
        \noisestate_0/dectime[11]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_68 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[32]  (.A(
        \top_code_0_dds_configdata[15] ), .B(\DDS_0/dds_state_0/N_569 )
        , .C(\DDS_0/dds_state_0/N_312 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[32] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[9]  (.D(
        \top_code_0_dds_configdata[8] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[9]_net_1 ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_0  (.A(\ADC_c[10] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_0 ));
    NOR2 \noisestate_0/sw_acq2_RNO_1  (.A(\noisestate_0/CS[3]_net_1 ), 
        .B(\noisestate_0/CS[4]_net_1 ), .Y(\noisestate_0/N_233 ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_47  (.A(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[11] ));
    DFN0C0 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[2] ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add )
        , .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[2] ));
    NOR3B \scalestate_0/necount_LE_M_RNIPTOI_0  (.A(scalestate_0_ne_le)
        , .B(\scalestate_0/CS[12]_net_1 ), .C(
        \scalestate_0/necount_LE_M_net_1 ), .Y(
        \scalestate_0/timecount_13_sqmuxa_0 ));
    NOR2A \top_code_0/un1_xa_2_0_a2  (.A(\top_code_0/N_336 ), .B(
        \top_code_0/N_159 ), .Y(\top_code_0/un1_xa_2 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_8  (.A(
        \timer_top_0/dataout[9] ), .B(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_8_Y ));
    NOR2B \scalestate_0/strippluse_RNO[3]  (.A(\scalestate_0/N_562 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[3]_net_1 ));
    NOR3B \top_code_0/plusedata_1_sqmuxa_0_a2  (.A(\xa_c[7] ), .B(
        \top_code_0/plusedata_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_139 ), .Y(\top_code_0/plusedata_1_sqmuxa ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n13 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i14_mux ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[9]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[9] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_9_inst ), .S(top_code_0_n_s_ctrl_1), 
        .Y(\Signal_Noise_Acq_0_dataout[9] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[4]  (.A(
        \s_acq_change_0/s_acqnum_5[4] ), .B(
        \s_acq_change_0_s_acqnum[4] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_74 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[11]  (.D(
        \top_code_0_state_1ms_data[11] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[11]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_20[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[2]_net_1 ), .B(
        \pd_pluse_top_0/count_6[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_2[0] ));
    DFN1 \s_acq_change_0/s_load  (.D(
        \s_acq_change_0/s_load_0_0_RNIEJ0I1_net_1 ), .CLK(GLA_net_1), 
        .Q(s_acq_change_0_s_load));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m45_0 ));
    MX2 \scanstate_0/timecount_1_RNO_0[15]  (.A(
        \scanstate_0/dectime[15]_net_1 ), .B(
        \scanstate_0/acqtime[15]_net_1 ), .S(\scanstate_0/CS[4]_net_1 )
        , .Y(\scanstate_0/N_73 ));
    DFN1 \DUMP_OFF_0/off_on_timer_0/count[3]  (.D(
        \DUMP_OFF_0/off_on_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/count_3[3] ));
    NOR2B \state_1ms_0/timecount_RNO_5[7]  (.A(
        \state_1ms_0/PLUSECYCLE[7]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[7] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/fAND2_8_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_9_net ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_40_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_41_i ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_5  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_4_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_0_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_4_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_5_Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m42  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_39 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_42 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_43 ));
    MX2B \plusestate_0/timecount_1_RNO[2]  (.A(\plusestate_0/N_73 ), 
        .B(\plusestate_0/N_247 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[2] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIM8594[3]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_1[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_0[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_16[0] ));
    DFN1E1 \top_code_0/noisedata[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[11] ));
    AOI1 \scalestate_0/necount_LE_M_RNIBQQD  (.A(
        \scalestate_0/necount_LE_M_net_1 ), .B(
        \scalestate_0/CS[15]_net_1 ), .C(
        \scalestate_0/timecount_16_sqmuxa_1 ), .Y(
        \scalestate_0/necount_LE_M_RNIBQQD_net_1 ));
    DFN1E1 \plusestate_0/PLUSETIME[15]  (.D(\top_code_0_plusedata[15] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[15]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m57  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_54 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_57 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_58 ));
    IOTRI_OR_EB \Q2Q7_pad/U0/U1  (.D(
        \PLUSE_0/qq_state_1/Q1Q8_Q2Q7_RNO_0_net_1 ), .E(VCC), .OCLK(
        GLA_net_1), .DOUT(\Q2Q7_pad/U0/NET1 ), .EOUT(
        \Q2Q7_pad/U0/NET2 ));
    AO1 \scalestate_0/timecount_ret_81_RNO  (.A(
        \scalestate_0/CUTTIME180[4]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[4] ), .Y(
        \scalestate_0/timecount_20_iv_2[4] ));
    NOR2B \scalestate_0/timecount_ret_59_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[0]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[0] ));
    MX2 \scalestate_0/s_acq_RNO_0  (.A(\scalestate_0/N_1197 ), .B(
        scalestate_0_s_acq), .S(\scalestate_0/N_1169 ), .Y(
        \scalestate_0/N_724 ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIFG5N[1]  (.A(
        \DUMP_0/count_1[1] ), .B(\DUMP_0/count_1[0] ), .Y(
        \DUMP_0/dump_timer_0/count_c1 ));
    MX2 \state1ms_choice_0/bri_cycle_RNO_0  (.A(PLUSE_0_bri_cycle), .B(
        state_1ms_0_bri_cycle), .S(top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/bri_cycle_5 ));
    OR2B \PLUSE_0/qq_state_0/cs_RNIB5QN[3]  (.A(\PLUSE_0/i_4[3] ), .B(
        \PLUSE_0/qq_state_0/cs[3]_net_1 ), .Y(
        \PLUSE_0/qq_state_0/N_79 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_4_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_89_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_87_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_4_inst ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m235  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_236 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[6]  (.A(
        \scanstate_0_timecount[6] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_211 ));
    NOR2B \DDS_0/dds_state_0/para_RNO_0[7]  (.A(
        \DDS_0/dds_state_0/para[8]_net_1 ), .B(
        \DDS_0/dds_state_0/N_534 ), .Y(\DDS_0/dds_state_0/N_273 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[6]  (.A(
        \state_1ms_0_timecount[6] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_212 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m211  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_208 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_211 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_212 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[16]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[16]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[6]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m257  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[15] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_258 ));
    NOR3C \scalestate_0/timecount_ret_22_RNO_0  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[10]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[10] ));
    MX2B \noisestate_0/rt_sw_RNO_0  (.A(noisestate_0_rt_sw), .B(
        \noisestate_0/CS[5]_net_1 ), .S(\noisestate_0/N_248 ), .Y(
        \noisestate_0/N_110 ));
    DFN1 \top_code_0/pluse_rst_0_0  (.D(
        \top_code_0/pluse_rst_0_0_RNIO7ND3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_pluse_rst_0));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[4]  (.A(
        \state_1ms_0_timecount[4] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_222 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[11] ));
    DFN1E1 \top_code_0/s_addchoice[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice[1] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[14]_net_1 ));
    DFN1 \PLUSE_0/qq_timer_0/count[1]  (.D(
        \PLUSE_0/qq_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_9[1] ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[3]  (.D(
        \DUMP_0/dump_coder_0/para4_4[3]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[3]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[6]  (.A(
        \noisestate_0/acqtime[6]_net_1 ), .B(
        \noisestate_0/dectime[6]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_63 ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[6]  (.D(
        \DUMP_0/dump_coder_0/para5_4[6] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[6]_net_1 ));
    OA1A \plusestate_0/tetw_pluse_RNO  (.A(\plusestate_0/N_302 ), .B(
        plusestate_0_tetw_pluse), .C(top_code_0_pluse_rst), .Y(
        \plusestate_0/tetw_pluse_RNO_0 ));
    AX1C \ClockManagement_0/clk_div500_0/un1_count_1_I_36  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_11[0] ), 
        .B(\ClockManagement_0/clk_div500_0/count[6]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/I_36 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[1]  (.D(
        \DUMP_0/dump_coder_0/para2_4[1]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[1]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO[18]  (.A(\state_1ms_0/N_85 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[18]_net_1 ));
    OR2B \top_code_0/un1_state_1ms_rst_n117_47_i_o2_0  (.A(\xa_c[3] ), 
        .B(\xa_c[1] ), .Y(\top_code_0/N_149 ));
    NOR2B \state_1ms_0/timecount_RNO_6[15]  (.A(
        \state_1ms_0/PLUSETIME[15]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[15] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_12  (.A(\xd_in[2] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[2] ));
    XOR2 \PLUSE_0/qq_coder_1/i_reg10_2[0]  (.A(\PLUSE_0/qq_para3[2] ), 
        .B(\PLUSE_0/count_7[2] ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_2[0]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m65  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_58 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_65 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_66 ));
    DFN1E1 \noisestate_0/dectime[12]  (.D(\top_code_0_noisedata[12] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[12]_net_1 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i2_mux ));
    DFN1E1 \scalestate_0/CUTTIME90[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[15]_net_1 ));
    OA1B \noisestate_0/CS_RNO[4]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[4]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[4] )
        , .Y(\noisestate_0/CS_RNO[4]_net_1 ));
    DFN1E1 \noisestate_0/timecount_1[10]  (.D(
        \noisestate_0/timecount_5[10] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[10] ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[0]  (
        .D(\top_code_0_s_periodnum[0] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[0]_net_1 )
        );
    NOR2A \DDS_0/dds_state_0/para_RNO_3[16]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[15] )
        , .Y(\DDS_0/dds_state_0/N_294 ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BFF1_1_inst  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ));
    IOTRI_OB_EB \relay_close_pad[5]/U0/U1  (.D(\relay_close_c[5] ), .E(
        VCC), .DOUT(\relay_close_pad[5]/U0/NET1 ), .EOUT(
        \relay_close_pad[5]/U0/NET2 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[15]  (.A(
        \timer_top_0/state_switch_0/N_187 ), .B(
        \timer_top_0/state_switch_0/N_189 ), .C(
        \timer_top_0/state_switch_0/N_188 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[15] ));
    MAJ3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I1_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[1]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[1] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I0_un1_CO1 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N142 ));
    NOR2B \DUMP_OFF_0/off_on_coder_0/i_RNO[0]  (.A(
        bri_dump_sw_0_dumpoff_ctr), .B(bri_dump_sw_0_reset_out), .Y(
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[0] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_26  (.A(
        \timer_top_0/dataout[20] ), .B(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_26_Y ));
    NOR3C \DUMP_0/dump_coder_0/para5_RNIFUGAG[0]  (.A(
        state1ms_choice_0_reset_out), .B(
        \DUMP_0/dump_coder_0/i_reg16_NE[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/N_19 ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_6  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/NE_NUM[9]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_6_Y ));
    DFN1 \scalestate_0/fst_lst_pulse  (.D(
        \scalestate_0/fst_lst_pulse_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/fst_lst_pulse_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[2] ));
    IOTRI_OB_EB \syn_md_tmp_pad/U0/U1  (.D(syn_md_tmp_c), .E(VCC), 
        .DOUT(\syn_md_tmp_pad/U0/NET1 ), .EOUT(
        \syn_md_tmp_pad/U0/NET2 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_33  (.A(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ));
    AO1B \state_1ms_0/CS_RNO_0[1]  (.A(\state_1ms_0/CS_i[0]_net_1 ), 
        .B(timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[1] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[18]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[18]_net_1 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[8]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[12]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[12]_net_1 ), .CLK(
        ddsclkout_c), .Q(
        \pd_pluse_top_0/pd_pluse_state_0/cs[12]_net_1 ));
    DFN1E1 \top_code_0/sigtimedata[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[12] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIFSMN7[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_12[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[8]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[8]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_284 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[19]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_56 ), .Y(
        \timer_top_0/timer_0/timedata_4[19] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_50_i ));
    DFN1E0 \DDS_0/dds_state_0/para[24]  (.D(\DDS_0/dds_state_0/N_23 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[24]_net_1 ));
    OR2A \state_1ms_0/timecount_RNO[0]  (.A(top_code_0_state_1ms_rst_n)
        , .B(\state_1ms_0/N_67 ), .Y(
        \state_1ms_0/timecount_RNO[0]_net_1 ));
    NOR2 \scalestate_0/CS_RNITQUB[4]  (.A(\scalestate_0/CS[4]_net_1 ), 
        .B(\scalestate_0/CS[10]_net_1 ), .Y(\scalestate_0/N_1263 ));
    XA1 \DUMP_OFF_0/off_on_timer_0/count_RNO[3]  (.A(
        \DUMP_OFF_0/off_on_timer_0/count_c2 ), .B(
        \DUMP_OFF_0/count_3[3] ), .C(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_n3 ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIEKJD1[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_0[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_1[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_8[0] ));
    XO1 \PLUSE_0/qq_coder_0/un1_qq_para2_NE_1[0]  (.A(
        \PLUSE_0/count_9[3] ), .B(\PLUSE_0/qq_para2[3] ), .C(
        \PLUSE_0/qq_coder_0/un1_qq_para2_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_1[0]_net_1 ));
    DFN1 \noisestate_0/CS[4]  (.D(\noisestate_0/CS_RNO[4]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[4]_net_1 ));
    DFN1E1 \scalestate_0/NE_NUM[3]  (.D(\top_code_0_scaledatain[3] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[3]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[6] ));
    MX2 \state_1ms_0/timecount_RNO_0[16]  (.A(
        \state_1ms_0/timecount_8[16] ), .B(\state_1ms_0_timecount[16] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_83 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[7]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[7]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_2[7] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[2]  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n2 ));
    DFN1E1 \top_code_0/halfdata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[6] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m25  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_24 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_25 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_26 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIUDTT[7]  (
        .A(\pd_pluse_top_0/count_1[7] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[7]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_5[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_3[0] ));
    AO1C \state_1ms_0/timecount_RNO_3[5]  (.A(
        \state_1ms_0/M_DUMPTIME[5]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_i[0]_net_1 ), 
        .Y(\state_1ms_0/timecount_8_iv_0[5] ));
    AO1A \scanstate_0/calctrl_RNO_0  (.A(\scanstate_0/CS[5]_net_1 ), 
        .B(scanstate_0_calctrl), .C(\scanstate_0/CS[2]_net_1 ), .Y(
        \scanstate_0/N_131 ));
    MX2A \pd_pluse_top_0/pd_pluse_state_0/en1_RNO_1  (.A(
        \pd_pluse_top_0/i_1[2] ), .B(\pd_pluse_top_0/i_1[3] ), .S(
        \pd_pluse_top_0/pd_pluse_state_0/N_166 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/en1_0_i_1 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]  (
        .D(\top_code_0_n_acqnum_2[11] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]_net_1 )
        );
    NOR3B \top_code_0/state_1ms_lc_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/state_1ms_lc_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_152 ), .Y(\top_code_0/state_1ms_lc_1_sqmuxa ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNIFLVR2[6]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c4 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c6 ));
    DFN1E1 \plusestate_0/DUMPTIME[3]  (.D(\top_code_0_plusedata[3] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[3]_net_1 ));
    DFN1 \scalestate_0/CS[3]  (.D(\scalestate_0/CS_RNO_1[3] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[3]_net_1 ));
    IOTRI_OB_EB \relay_on_pad[1]/U0/U1  (.D(\relay_on_c[1] ), .E(VCC), 
        .DOUT(\relay_on_pad[1]/U0/NET1 ), .EOUT(
        \relay_on_pad[1]/U0/NET2 ));
    MX2 \plusestate_0/timecount_1_RNO_0[7]  (.A(
        \plusestate_0/DUMPTIME[7]_net_1 ), .B(
        \plusestate_0/PLUSETIME[7]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_78 ));
    OR3 \DUMP_0/dump_coder_0/para6_RNIGKPR2[0]  (.A(
        \DUMP_0/dump_coder_0/i_reg16_10[0] ), .B(
        \DUMP_0/dump_coder_0/i_reg16_0[0] ), .C(
        \DUMP_0/dump_coder_0/i_reg16_NE_5[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_8[0] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[15]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i20_mux ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_10_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_10_net ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[4]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_31_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[4] ));
    AND2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_35  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[1]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[2] ));
    DFN1E1 \top_code_0/noisedata[14]  (.D(\GPMI_0_dataout[14] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[14] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[9] ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[5]  (
        .D(\s_acq_change_0_s_acqnum[5] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[5]_net_1 )
        );
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_39  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[2]_net_1 ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[5] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[6] ));
    AO1 \scalestate_0/timecount_ret_73_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[7]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[7] ), .Y(
        \scalestate_0/timecount_20_iv_4[7] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_14[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[4]_net_1 ), .B(
        \pd_pluse_top_0/count_6[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_4[0] ));
    DFN1 \timer_top_0/state_switch_0/state_start  (.D(
        \timer_top_0/state_switch_0/state_start5 ), .CLK(GLA_net_1), 
        .Q(\timer_top_0/state_switch_0_state_start ));
    MX2A \state_1ms_0/timecount_RNO_0[5]  (.A(
        \state_1ms_0/timecount_8_iv[5] ), .B(
        \state_1ms_0_timecount[5] ), .S(\state_1ms_0/CS[9]_net_1 ), .Y(
        \state_1ms_0/N_72 ));
    DFN1E1 \top_code_0/noisedata[13]  (.D(\GPMI_0_dataout[13] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[13] ));
    DFN1 \state1ms_choice_0/pluse_start  (.D(
        \state1ms_choice_0/pluse_start_RNO_1 ), .CLK(GLA_net_1), .Q(
        bri_div_start_0));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_11_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_14_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_11_net ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI2B5C[1]  
        (.A(\s_acq_change_0_s_stripnum[0] ), .B(
        \s_acq_change_0_s_stripnum[1] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_1 ));
    NOR2A \scanstate_0/CS_RNI97DM_0[1]  (.A(net_33), .B(
        \scanstate_0/CS[1]_net_1 ), .Y(\scanstate_0/timecount_cnst[2] )
        );
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m47_2 ));
    NOR2B \DDS_0/dds_coder_0/i_RNO[0]  (.A(dds_change_0_dds_conf), .B(
        dds_change_0_dds_rst), .Y(\DDS_0/dds_coder_0/i_RNO[0]_net_1 ));
    NOR3A \syn_md_module_1/syn_md_0/count_RNIV9NM[3]  (.A(
        \syn_md_module_1/syn_md_0/N_52 ), .B(
        \syn_md_module_1/syn_md_0/N_18 ), .C(
        \syn_md_module_1/syn_md_0/count[3]_net_1 ), .Y(
        \syn_md_module_1/syn_md_0/N_50 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m42 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[9]_net_1 ));
    NOR2B \ClockManagement_0/clk_div500_0/count_RNINJ1O[7]  (.A(
        \ClockManagement_0/clk_div500_0/count[6]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_2 ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_11[10]  (.A(
        \sd_acq_top_0/count_0[12] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[12]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_7[10] ));
    DFN1 \DUMP_0/dump_timer_0/count[8]  (.D(
        \DUMP_0/dump_timer_0/count_n8 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count[8] ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[7]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[7] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_7_inst ), .S(top_code_0_n_s_ctrl_1), 
        .Y(\Signal_Noise_Acq_0_dataout[7] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[12]  (.A(
        \timer_top_0/state_switch_0/N_257 ), .B(
        \timer_top_0/state_switch_0/N_259 ), .C(
        \timer_top_0/state_switch_0/N_258 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[12] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[7]  (.A(
        \scalestate_0_strippluse[7] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[7] ));
    NOR3C \scalestate_0/timecount_20_iv_5_RNO_1[4]  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[4]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[4] ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[5]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[5] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[5] ));
    NOR3 \scalestate_0/necount_cmp_0/NOR3_0  (.A(
        \scalestate_0/necount_cmp_0/OA1A_0_Y ), .B(
        \scalestate_0/necount_cmp_0/AND2A_0_Y ), .C(
        \scalestate_0/necount_cmp_0/OA1C_0_Y ), .Y(
        \scalestate_0/necount_cmp_0/NOR3_0_Y ));
    DFN1 \DUMP_0/dump_timer_0/count[1]  (.D(
        \DUMP_0/dump_timer_0/count_n1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_1[1] ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/count[3]  (.D(
        \DSTimer_0/dump_sustain_timer_0/count_n3 ), .CLK(clock_10khz), 
        .Q(\DSTimer_0/dump_sustain_timer_0/count[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n11 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11]/Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m255  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_254 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_255 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_256 ));
    AO1 \DDS_0/dds_state_0/para_RNO[34]  (.A(
        \DDS_0/dds_state_0/para[34]_net_1 ), .B(
        \DDS_0/dds_state_0/N_538_0 ), .C(\DDS_0/dds_state_0/N_524 ), 
        .Y(\DDS_0/dds_state_0/para_9[34] ));
    OA1 \scanstate_0/s_acq_RNO  (.A(\scanstate_0/CS[4]_net_1 ), .B(
        scanstate_0_s_acq), .C(net_33_0), .Y(\scanstate_0/s_acq_RNO_0 )
        );
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[20]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[20]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n8 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8]/Y ));
    AX1C \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_3_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/count_10[3] ), .C(\sd_acq_top_0/count_10[4] ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/count1[4] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_0  (.A(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .B(
        \timer_top_0/dataout[5] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_0_Y ));
    NOR2B \state_1ms_0/timecount_RNO_6[3]  (.A(
        \state_1ms_0/CUTTIME[3]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[3] ));
    AO1B \state_1ms_0/timecount_RNO_3[3]  (.A(
        \state_1ms_0/M_DUMPTIME[3]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_i[0]_net_1 ), 
        .Y(\state_1ms_0/timecount_8_iv_0[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[7] ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[20]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[20] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[20] ));
    DFN1 \scanstate_0/s_acq  (.D(\scanstate_0/s_acq_RNO_0 ), .CLK(
        GLA_net_1), .Q(scanstate_0_s_acq));
    NOR2 \top_code_0/un1_xa_8_16_i_i_o3_i_a2_1  (.A(\xa_c[17] ), .B(
        \xa_c[16] ), .Y(\top_code_0/un1_xa_8_16_i_i_o3_i_a2_1_net_1 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[15]  (.A(
        \s_acq_change_0/s_acqnum_5[15] ), .B(
        \s_acq_change_0_s_acqnum[15] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_85 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_9  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[2] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m202  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_201 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_202 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_203 ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNIS6241[8]  (.A(
        \ClockManagement_0/clk_div500_0/count[2]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[8]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count[3]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_4 ));
    NOR2B \DDS_0/dds_state_0/para_RNO[36]  (.A(
        \DDS_0/dds_state_0/para[36]_net_1 ), .B(
        \DDS_0/dds_state_0/N_538_1 ), .Y(
        \DDS_0/dds_state_0/para_9[36] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m70  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_69 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_70 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_71 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[16]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[16]_net_1 ));
    NOR3B \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[8]  (.A(
        \pd_pluse_top_0/i_0[5] ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_i[0]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[8] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIMF1G[1]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[1]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_0[0] ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_3  (.A(\ADC_c[7] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_3 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[10]  (.A(
        \top_code_0_s_acqnum_2[10] ), .B(\scalestate_0_s_acqnum[10] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[10] ));
    NOR2B \plusestate_0/DUMPTIME_1_sqmuxa  (.A(top_code_0_pluse_lc), 
        .B(top_code_0_pluseload), .Y(
        \plusestate_0/DUMPTIME_1_sqmuxa_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m42 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[17] ));
    DFN1E1 \scanstate_0/acqtime[0]  (.D(\top_code_0_scandata[0] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[0]_net_1 ));
    AO1A \topctrlchange_0/sw_acq2_RNO_1  (.A(scalestate_0_sw_acq2), .B(
        \top_code_0_change_0[0] ), .C(\topctrlchange_0/sw_acq2in1_i_m )
        , .Y(\topctrlchange_0/sw_acq2_6_iv ));
    NOR2 \top_code_0/scan_start_ret_3_RNO_0  (.A(\top_code_0/N_144 ), 
        .B(\top_code_0/N_149 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_47_i_a2_0 ));
    NOR3A \top_code_0/dump_sustain_data_1_sqmuxa_0_a2  (.A(
        \top_code_0/cal_data_1_sqmuxa_1 ), .B(\top_code_0/N_144 ), .C(
        \top_code_0/N_167 ), .Y(
        \top_code_0/dump_sustain_data_1_sqmuxa ));
    XA1C \PLUSE_0/qq_coder_0/i_RNO_1[1]  (.A(\PLUSE_0/count_9[2] ), .B(
        \PLUSE_0/qq_para1[2] ), .C(\PLUSE_0/qq_coder_0/un1_count_1[0] )
        , .Y(\PLUSE_0/qq_coder_0/i_0_1[1] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[7]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO[20]  (.A(
        \scalestate_0_timecount[20] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[20]_net_1 ));
    MX2 \scalestate_0/necount_RNO_0[4]  (.A(\scalestate_0/necount1[4] )
        , .B(\scalestate_0/necount[4]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_734 ));
    MX2 \plusestate_0/timecount_1_RNO_0[9]  (.A(
        \plusestate_0/PLUSETIME[9]_net_1 ), .B(
        \plusestate_0/DUMPTIME[9]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_80 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m47 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[6]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[6]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/en2 ));
    IOPAD_TRI \dumpoff_pad/U0/U0  (.D(\dumpoff_pad/U0/NET1 ), .E(
        \dumpoff_pad/U0/NET2 ), .PAD(dumpoff));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_38_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m44_3 ));
    NOR2 \DUMP_ON_0/off_on_coder_0/i_RNO_1[1]  (.A(
        \DUMP_ON_0/count_5[1] ), .B(\DUMP_ON_0/count_5[0] ), .Y(
        \DUMP_ON_0/off_on_coder_0/i_0_1[1] ));
    OR3 \dds_change_0/dds_rst_RNO_1  (.A(\dds_change_0/ddsrstin2_m ), 
        .B(\dds_change_0/ddsrstin3_m ), .C(\dds_change_0/ddsrstin1_m ), 
        .Y(\dds_change_0/dds_rst_6 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m220  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_221 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNICUCH[17]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[17]_net_1 ), .B(
        \sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_17[0] ));
    NOR2B \scalestate_0/necount_LE_M_RNI1CBP  (.A(
        \scalestate_0/timecount_12_sqmuxa_0 ), .B(
        top_code_0_scale_rst_0), .Y(\scalestate_0/N_258_0 ));
    DFN1E1 \scalestate_0/M_NUM[4]  (.D(\top_code_0_scaledatain[4] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[4]_net_1 ));
    NOR2B \CAL_0/cal_div_0/cal_RNO  (.A(\CAL_0/cal_div_0/N_35 ), .B(
        net_33), .Y(\CAL_0/cal_div_0/cal_RNO_net_1 ));
    NOR3 \top_code_0/state_1ms_load_RNO_1  (.A(\top_code_0/N_152 ), .B(
        \top_code_0/N_163 ), .C(\top_code_0/N_147 ), .Y(
        \top_code_0/N_314 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_3_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_3_net ));
    OR2A \top_code_0/sd_sacq_choice_1_sqmuxa_0_o2  (.A(\xa_c[4] ), .B(
        \top_code_0/N_142 ), .Y(\top_code_0/N_163 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m54  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_55 ));
    NOR2A \scalestate_0/timecount_ret_73_RNO_4  (.A(
        \scalestate_0/CUTTIME90[7]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[7] ));
    OR3 \state_1ms_0/timecount_RNO_1[3]  (.A(
        \state_1ms_0/timecount_8_iv_1[3] ), .B(
        \state_1ms_0/timecount_8_iv_0[3] ), .C(
        \state_1ms_0/timecount_8_iv_2[3] ), .Y(
        \state_1ms_0/timecount_8[3] ));
    DFN1 \ClockManagement_0/clk_div500_0/count[6]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[6] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[6]_net_1 ));
    DFN1E1 \top_code_0/halfdata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[5] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_34  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[7] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[6] )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2 ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_70_i ));
    NOR2B \scalestate_0/timecount_ret_65_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[13]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[13] ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        );
    OR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[9]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .B(
        \sd_acq_top_0/i_5[2] ), .C(\sd_acq_top_0/i_5[3] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_207 ));
    NOR2B \state_1ms_0/timecount_RNO[8]  (.A(\state_1ms_0/N_75 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[8]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[8] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_62_i ));
    AND3 \scalestate_0/necount_cmp_1/AND3_1  (.A(
        \scalestate_0/necount_cmp_1/XNOR2_8_Y ), .B(
        \scalestate_0/necount_cmp_1/XNOR2_5_Y ), .C(
        \scalestate_0/necount_cmp_1/XNOR2_3_Y ), .Y(
        \scalestate_0/necount_cmp_1/AND3_1_Y ));
    OR3B \scalestate_0/fst_lst_pulse_RNIR20M2  (.A(
        timer_top_0_clk_en_scale_0), .B(\scalestate_0/N_1309 ), .C(
        \scalestate_0/sw_acq1_1_sqmuxa ), .Y(\scalestate_0/un1_CS6_34 )
        );
    DFN1E0 \DDS_0/dds_state_0/para[33]  (.D(
        \DDS_0/dds_state_0/para_9[33] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[33]_net_1 ));
    AOI1B \PLUSE_0/qq_state_0/cs_RNO[1]  (.A(
        \PLUSE_0/qq_state_0/cs_i[0]_net_1 ), .B(
        \PLUSE_0/qq_state_0/N_82 ), .C(\PLUSE_0/qq_state_0/cs4 ), .Y(
        \PLUSE_0/qq_state_0/cs_RNO_1[1] ));
    DFN1 \plusestate_0/pluse_acq  (.D(
        \plusestate_0/pluse_acq_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        plusestate_0_pluse_acq));
    DFN1E0 \DUMP_0/dump_coder_0/para2[11]  (.D(
        \DUMP_0/dump_coder_0/para2_4[11]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[11]_net_1 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_14  (.A(
        \timer_top_0/dataout[18] ), .B(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_14_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m44_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[15] ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_23[10]  (.A(
        \sd_acq_top_0/count_1[9] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[9]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_3[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_10[10] ));
    IOTRI_OB_EB \sigtimeup_pad/U0/U1  (.D(sigtimeup_c), .E(VCC), .DOUT(
        \sigtimeup_pad/U0/NET1 ), .EOUT(\sigtimeup_pad/U0/NET2 ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_11_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_14_net ), 
        .B(\pd_pluse_top_0/count[14] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[14] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i18_mux ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIQT421[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_2[0] ));
    NOR2A \scalestate_0/timecount_ret_29_RNO_4  (.A(
        \scalestate_0/CUTTIME90[1]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[1] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m123  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[19] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_124 ));
    NOR3C \scalestate_0/timecount_ret_57_RNO_3  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[0]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[0] ));
    NOR2A \timer_top_0/state_switch_0/state_over_n_RNO_1  (.A(
        \timer_top_0/state_switch_0/N_295 ), .B(
        scanstate_0_state_over_n), .Y(
        \timer_top_0/state_switch_0/N_279 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[0]  (.A(
        \timer_top_0/state_switch_0/N_242 ), .B(
        \timer_top_0/state_switch_0/N_244 ), .C(
        \timer_top_0/state_switch_0/N_243 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[0] ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_52_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[1] )
        );
    MX2 \scalestate_0/s_acqnum_1_RNO_1[0]  (.A(\scalestate_0/N_448 ), 
        .B(\scalestate_0/ACQECHO_NUM[0]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[0] ));
    DFN1 \scalestate_0/intertodsp  (.D(
        \scalestate_0/intertodsp_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        calcuinter_c));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[1]  (.A(
        \scalestate_0_strippluse[1] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[1] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_113  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_12_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_144_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_113_Y ));
    NOR3C \scalestate_0/timecount_ret_56_RNO_1  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[19]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[19] ));
    NOR2 \plusestate_0/CS_RNIN1IP[6]  (.A(\plusestate_0/CS[7]_net_1 ), 
        .B(\plusestate_0/CS[6]_net_1 ), .Y(\plusestate_0/N_302 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[10] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i6_mux ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[28]  (.D(
        \top_code_0_dds_configdata[11] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[28]_net_1 ));
    NOR2B \scalestate_0/CS_RNO[19]  (.A(\scalestate_0/N_1231 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[19]_net_1 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[15]  (.A(
        \timer_top_0/state_switch_0/N_185 ), .B(
        \timer_top_0/state_switch_0/N_186 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[15] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[15]_net_1 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m47_5 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_61  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_55_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_43_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_61_Y ));
    OR3 \scalestate_0/timecount_ret_53_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[18] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[18] ), .C(
        \scalestate_0/timecount_20_0_iv_2[18] ), .Y(
        \scalestate_0/timecount_20_0_iv_4[18] ));
    DFN1E1 \top_code_0/plusedata[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[11] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[4]  (.D(
        \top_code_0_n_divnum_0[4] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[4]_net_1 ));
    DFN1 \DDS_0/dds_timer_0/count[5]  (.D(\DDS_0/dds_timer_0/count_n5 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[5] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/entop_RNO  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/entop_RNO_net_1 )
        );
    NOR2A \scalestate_0/strippluse_RNO_1[9]  (.A(\scalestate_0/N_429 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[9] ));
    DFN1E1 \top_code_0/s_acqnum[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[0] ));
    NOR2A \scalestate_0/timecount_ret_62_RNO_4  (.A(
        \scalestate_0/CUTTIME90[12]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[12] ));
    NOR2B \nsctrl_choice_0/dumpoff_ctr_RNO  (.A(
        \nsctrl_choice_0/dumpoff_ctr_5 ), .B(net_27), .Y(
        \nsctrl_choice_0/dumpoff_ctr_RNO_1 ));
    OR2B \DDS_0/dds_state_0/cs_RNO_0[2]  (.A(\DDS_0/i[1] ), .B(
        \DDS_0/dds_state_0/cs[1]_net_1 ), .Y(\DDS_0/dds_state_0/N_228 )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI8QCH[15]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[15]_net_1 ), .B(
        \sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_15[0] ));
    DFN1E1 \scalestate_0/CUTTIME90[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[10]_net_1 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[15]  (.D(
        \top_code_0_state_1ms_data[15] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[15]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/stateover  (.D(
        \sd_acq_top_0/sd_sacq_state_0/stateover_RNO_2 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/sd_sacq_state_0_stateover ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[1] ));
    DFN1E1 \scanstate_0/timecount_1[14]  (.D(
        \scanstate_0/timecount_5[14] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[14] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[2]  (.A(
        \scalestate_0/ACQ180_NUM[2]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[2]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_450 ));
    OR3 \scalestate_0/timecount_ret_79_RNO  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_6_0 ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_6_1 ), .C(
        \scalestate_0/un1_timecount_2_sqmuxa_7 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_9 ));
    XA1 \DUMP_OFF_1/off_on_timer_0/count_RNO[2]  (.A(
        \DUMP_OFF_1/off_on_timer_0/count_c1 ), .B(
        \DUMP_OFF_1/count_4[2] ), .C(
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_n2 ));
    DFN1E1 \top_code_0/plusedata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[5] ));
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_5  (.A(
        \scalestate_0/NE_NUM[1]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .C(
        \scalestate_0/necount_cmp_1/OR2A_1_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_5_Y ));
    IOPAD_TRI \relay_close_pad[0]/U0/U0  (.D(
        \relay_close_pad[0]/U0/NET1 ), .E(\relay_close_pad[0]/U0/NET2 )
        , .PAD(relay_close[0]));
    MAJ3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I2_un1_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[2]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[2] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N142 ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I2_un1_CO1 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_7[3]  (.A(
        \DUMP_0/dump_coder_0/para1[2]_net_1 ), .B(\DUMP_0/count_1[2] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_2[0] ));
    NOR2A \DUMP_0/dump_coder_0/i_RNO[6]  (.A(
        \DUMP_0/dump_coder_0/N_19 ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO[6]_net_1 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[11]  (.A(
        \DDS_0/dds_state_0/N_328 ), .B(\DDS_0/dds_state_0/N_327 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[11] ), .Y(
        \DDS_0/dds_state_0/N_87 ));
    NOR2B \PLUSE_0/qq_timer_1/count_RNI8L8E1[2]  (.A(
        \PLUSE_0/qq_timer_1/count_c1 ), .B(\PLUSE_0/count_7[2] ), .Y(
        \PLUSE_0/qq_timer_1/count_c2 ));
    NOR2A \DUMP_0/dump_coder_0/i_RNO_0[4]  (.A(
        \DUMP_0/dump_coder_0/un1_count_2_NE[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_3_i[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_0[4] ));
    AND3 \scalestate_0/necount_cmp_1/AND3_2  (.A(
        \scalestate_0/necount_cmp_1/XNOR2_0_Y ), .B(
        \scalestate_0/necount_cmp_1/XNOR2_9_Y ), .C(
        \scalestate_0/necount_cmp_1/XNOR2_7_Y ), .Y(
        \scalestate_0/necount_cmp_1/AND3_2_Y ));
    DFN1E1 \scalestate_0/CUTTIME180[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[15]_net_1 )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i22_mux ));
    NOR2B \DDS_0/dds_coder_0/m12_0  (.A(\DDS_0/count[1] ), .B(
        \DDS_0/count[3] ), .Y(\DDS_0/dds_coder_0/m12_0_net_1 ));
    OR3 \bridge_div_0/count_RNIRP683[3]  (.A(
        \bridge_div_0/clear1_n17_NE_0[0] ), .B(
        \bridge_div_0/clear1_n17_0[0] ), .C(
        \bridge_div_0/clear1_n17_NE_1[0] ), .Y(
        \bridge_div_0/clear1_n17_NE[0] ));
    NOR3B \state_1ms_0/M_DUMPTIME_1_sqmuxa_0_a2  (.A(
        \top_code_0_state_1ms_lc[1] ), .B(\state_1ms_0/N_17 ), .C(
        \top_code_0_state_1ms_lc[0] ), .Y(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ));
    OR2A \scalestate_0/CS_RNIR4SG_0[12]  (.A(
        \scalestate_0/CS[12]_net_1 ), .B(scalestate_0_ne_le), .Y(
        \scalestate_0/N_1208 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[11]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[11] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_0[11] ));
    AO1A \state_1ms_0/timecount_RNO_2[2]  (.A(
        \state_1ms_0/PLUSECYCLE[2]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/PLUSETIME_i_m[2] ), 
        .Y(\state_1ms_0/timecount_8_iv_1[2] ));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_31  (.A(
        \ClockManagement_0/clk_10k_0/count[4]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] ), .Y(
        \ClockManagement_0/clk_10k_0/I_31_0 ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[2]  (.A(\i_6[1] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[2]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_215 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m282  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_281 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_282 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_283 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[15]  
        (.D(\s_acq_change_0_s_acqnum[15] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[15]_net_1 )
        );
    NOR3C \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_2_i ));
    NOR3C \PLUSE_0/qq_timer_0/count_0_sqmuxa  (.A(
        \PLUSE_0/qq_state_0_stateover ), .B(\PLUSE_0/up ), .C(
        bri_dump_sw_0_reset_out_0), .Y(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m78  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_79 ));
    DFN1 \ClockManagement_0/clk_10k_0/clk_5M_reg1  (.D(
        \ClockManagement_0/clk_10k_0/clk_5M_reg1_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(\ClockManagement_0/clk_10k_0/clk_5M_reg1_net_1 )
        );
    DFN1E1 \top_code_0/s_addchoice_1[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_1[0] ));
    OR2 \top_code_0/s_addchoice_1_sqmuxa_0_o2  (.A(\xa_c[4] ), .B(
        \xa_c[2] ), .Y(\top_code_0/N_144 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[4]  (.A(
        \DDS_0/dds_state_0/para[4]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_315 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[4] ));
    DFN1E1 \top_code_0/n_acqnum[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[3] ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1_RNO_0  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I4_un1_CO1 ), 
        .B(\s_acq_change_0_s_stripnum[5] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_5 ));
    DFN1E1 \noisestate_0/timecount_1[12]  (.D(
        \noisestate_0/timecount_5[12] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[12] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_17  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_17_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI8BQ6[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[8]_net_1 ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_8[0] ));
    DFN1 \scalestate_0/long_opentime  (.D(
        \scalestate_0/long_opentime_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_long_opentime));
    DFN1E1 \top_code_0/scalechoice[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0[4] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[2]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[2] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_15_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_15_net ));
    DFN1P0 \syn_md_module_1/syn_md_edge_detect_0/sig_r1  (.D(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_i ), .CLK(
        GLA_net_1), .PRE(top_code_0_scale_rst_0), .Q(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r1_i_0 ));
    DFN1 \PLUSE_0/qq_timer_1/count[2]  (.D(
        \PLUSE_0/qq_timer_1/count_n2 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_7[2] ));
    DFN1E1 \top_code_0/dds_choice  (.D(\top_code_0/N_66 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_dds_choice));
    DFN1E1 \scalestate_0/timecount_ret_27  (.D(
        \scalestate_0/timecount_m3_e_1 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_m3_e_1_reto ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[21]  (.A(
        \top_code_0_dds_configdata[4] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_510 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[21] ));
    DFN1 \scalestate_0/off_test  (.D(
        \scalestate_0/off_test_RNO_1_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_off_test));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n6 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6]/Y ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[6]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[6] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_66_i ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[1]  (.D(
        \top_code_0_state_1ms_data[1] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[1]_net_1 ));
    AO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[1] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[0] )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_65 ));
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_1  (.A(
        \scalestate_0/necount_cmp_1/NOR3A_1_Y ), .B(
        \scalestate_0/necount_cmp_1/OR2A_3_Y ), .C(
        \scalestate_0/necount_cmp_1/NAND3A_3_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_1_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_12  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_12_Y ));
    DFN1 \scalestate_0/s_acqnum_1[6]  (.D(
        \scalestate_0/s_acqnum_1_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[6] ));
    NOR2A \top_code_0/un1_state_1ms_rst_n117_2_i_a2_3  (.A(
        GPMI_0_code_en), .B(\xa_c[6] ), .Y(\top_code_0/N_11_3 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m42_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[17] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i12_mux ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m112  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_105 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_112 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[4] ));
    NOR3A \sd_acq_top_0/sd_sacq_coder_0/i_RNO[9]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_i[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[9]_net_1 ));
    DFN1E1 \scanstate_0/acqtime[5]  (.D(\top_code_0_scandata[5] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[5]_net_1 ));
    DFN1E1 \top_code_0/n_acqnum[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[9] ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_33  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[7] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[8] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[10] )
        );
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7_116_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[2]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIUMEH[14]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[14]_net_1 )
        , .B(\pd_pluse_top_0/count[14] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_14[0] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[11]  (.A(
        \s_acq_change_0/N_67 ), .B(net_27), .Y(
        \s_acq_change_0/s_stripnum_RNO[11]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_52_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_96  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_96_Y ));
    NOR2B \PLUSE_0/qq_timer_0/count_RNI5QRU[2]  (.A(
        \PLUSE_0/qq_timer_0/count_c1 ), .B(\PLUSE_0/count_9[2] ), .Y(
        \PLUSE_0/qq_timer_0/count_c2 ));
    DFN1 \plusestate_0/CS[6]  (.D(\plusestate_0/CS_RNO_0[6]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[6]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_RNO[4]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_12_1 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[4] ));
    XA1B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_55  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[0]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4_0 ));
    DFN1E1 \top_code_0/scandata[12]  (.D(\GPMI_0_dataout[12] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[12] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m47_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_162  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_22_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_111_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_162_Y ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_58_i ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6_RNO  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N152 ), 
        .B(\s_acq_change_0_s_stripnum[6] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_6 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_53  (.A(
        \timer_top_0/timer_0/N_5 ), .B(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .Y(
        \timer_top_0/timer_0/I_53 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[17]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[17] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[17] ));
    DFN1E1 \plusestate_0/DUMPTIME[15]  (.D(\top_code_0_plusedata[15] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[15]_net_1 ));
    NOR3A \ClockManagement_0/clk_10k_0/count_RNIM27A1[8]  (.A(
        \ClockManagement_0/clk_10k_0/count[1]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[8]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/count[2]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_4 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m42_6 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[11]_net_1 ));
    MX2 \bri_dump_sw_0/phase_ctr_RNO_0  (.A(top_code_0_pn_change), .B(
        scalestate_0_pn_out), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/phase_ctr_5 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_0_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_0_net ));
    IOTRI_OB_EB \sw_acq1_pad/U0/U1  (.D(sw_acq1_c), .E(VCC), .DOUT(
        \sw_acq1_pad/U0/NET1 ), .EOUT(\sw_acq1_pad/U0/NET2 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[11] ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_1[0]  (.A(
        \sd_acq_top_0/count[20] ), .B(\sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_1[0]_net_1 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[9]  (.D(
        \top_code_0_state_1ms_data[9] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[9]_net_1 ));
    NOR2B \top_code_0/relay_close_RNO[3]  (.A(\top_code_0/N_822 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[3]_net_1 ));
    OA1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_16  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]_net_1 )
        , .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_3 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_7 ));
    OR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIDL47Q[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6 ));
    DFN1E1 \top_code_0/bri_datain[13]  (.D(\GPMI_0_dataout[13] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[13] ));
    DFN1E1 \top_code_0/scandata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[6] ));
    DFN1E1 \top_code_0/dds_configdata[7]  (.D(\GPMI_0_dataout[7] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[7] ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[4]  (.D(
        \DUMP_0/dump_coder_0/para4_4[4]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[4]_net_1 ));
    AO1A \scalestate_0/timecount_ret_72_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/S_DUMPTIME[7]_net_1 ), .C(
        \scalestate_0/timecount_20_iv_1[7] ), .Y(
        \scalestate_0/timecount_20_iv_6[7] ));
    DFN1E1 \scalestate_0/timecount_ret_13  (.D(
        \scalestate_0/timecount_cnst_m_0[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_cnst_m_0_reto[9] ));
    DFN1 \nsctrl_choice_0/intertodsp  (.D(
        \nsctrl_choice_0/intertodsp_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_intertodsp));
    AND2 \bridge_div_0/dataall_1_I_1  (.A(\top_code_0_scaleddsdiv[0] ), 
        .B(\top_code_0_scaleddsdiv[3] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_TMP[0] ));
    OR3 \DUMP_0/dump_coder_0/para5_RNIS1NE2[2]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_0[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_4_0[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE_3[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_7[0] ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNILJ563[1]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_2 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_4 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_9 ));
    AO1B \scanstate_0/state_over_n_RNO  (.A(scanstate_0_state_over_n), 
        .B(\scanstate_0/N_255 ), .C(net_33), .Y(
        \scanstate_0/state_over_n_RNO_1 ));
    DFN1E1 \scanstate_0/acqtime[9]  (.D(\top_code_0_scandata[9] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[9]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_145  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_4_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_104_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_145_Y ));
    XA1C \DUMP_0/dump_coder_0/i_RNO_11[3]  (.A(\DUMP_0/count_0[7] ), 
        .B(\DUMP_0/dump_coder_0/para1[7]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_6[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_5[3] ));
    OR3 \state_1ms_0/timecount_RNO_1[11]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[11] ), .B(
        \state_1ms_0/CUTTIME_m[11] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[11] ), .Y(
        \state_1ms_0/timecount_8[11] ));
    DFN1E1 \top_code_0/n_acqnum[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[1] ));
    DFN1E1 \scalestate_0/timecount_ret_84  (.D(
        \scalestate_0/timecount_20_iv_2[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_2_reto[11] ));
    DFN1E0 \DDS_0/dds_state_0/para[4]  (.D(\DDS_0/dds_state_0/N_54 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[4]_net_1 ));
    DFN1 \DUMP_0/off_on_coder_1/i[0]  (.D(
        \DUMP_0/off_on_coder_1/i_RNO_1[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_1[0] ));
    MX2 \scalestate_0/CS_RNO_0[5]  (.A(\scalestate_0/CS[5]_net_1 ), .B(
        \scalestate_0/CS[4]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1220 ));
    IOTRI_OB_EB \relay_close_pad[1]/U0/U1  (.D(\relay_close_c[1] ), .E(
        VCC), .DOUT(\relay_close_pad[1]/U0/NET1 ), .EOUT(
        \relay_close_pad[1]/U0/NET2 ));
    NOR3A \timer_top_0/state_switch_0/state_start5_0_0_a2_4  (.A(
        net_27), .B(top_code_0_pluse_str), .C(
        top_code_0_state_1ms_start), .Y(
        \timer_top_0/state_switch_0/N_284 ));
    DFN1E1 \scalestate_0/timecount_ret_22  (.D(
        \scalestate_0/timecount_20_iv_3[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_3_reto[10] ));
    NOR2B \scalestate_0/soft_d_RNO  (.A(\scalestate_0/N_543 ), .B(
        top_code_0_scale_rst_3), .Y(\scalestate_0/soft_d_RNO_2 ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[9]  (.A(
        \top_code_0_dumpdata_0[9] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[9]_net_1 ));
    AO1 \scalestate_0/timecount_ret_77_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[6]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[6] ), .Y(
        \scalestate_0/timecount_20_iv_4[6] ));
    NOR3 \top_code_0/dds_load_RNO_1  (.A(\top_code_0/N_142 ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_157 ), .Y(
        \top_code_0/N_276 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m40  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[0] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_41 ));
    NOR2 \top_code_0/un1_state_1ms_rst_n117_43_i_a3_0_0  (.A(\xa_c[3] )
        , .B(\top_code_0/N_140 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_43_i_a3_0_0_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_154  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_158_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_9_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_154_Y ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[9]  (.A(
        \timer_top_0/state_switch_0/N_202 ), .B(
        \timer_top_0/state_switch_0/N_204 ), .C(
        \timer_top_0/state_switch_0/N_203 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[9] ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[6]  (.D(
        \DUMP_0/dump_coder_0/para4_4[6]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[6]_net_1 ));
    DFN1E1 \top_code_0/n_acqnum[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[5] ));
    DFN1 \top_code_0/scan_start_ret  (.D(top_code_0_scan_start), .CLK(
        GLA_net_1), .Q(\top_code_0/top_code_0_scan_start_reto ));
    DFN1E1 \scalestate_0/S_DUMPTIME[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[0]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[8] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[13]  (.D(
        \top_code_0_pd_pluse_data[13] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[13]_net_1 ));
    AO1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_62_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4_0 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6_0 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[4]_net_1 ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIIR0R2[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_2[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_3[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_9[0] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[5] )
        );
    DFN1E1 \top_code_0/scandata[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[2] ));
    DFN1E1 \top_code_0/state_1ms_lc[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/state_1ms_lc_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_lc[3] ));
    DFN1E1 \scalestate_0/NE_NUM[6]  (.D(\top_code_0_scaledatain[6] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[6]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[23]  (.A(
        \top_code_0_dds_configdata[6] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_299 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[23] ));
    OR2A \top_code_0/un1_xa_2_0_o2  (.A(\xa_c[5] ), .B(\xa_c[7] ), .Y(
        \top_code_0/N_140 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNI4KTT[9]  (
        .A(\pd_pluse_top_0/count_0[9] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[9]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_6[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_5[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[6]_net_1 ));
    NOR2B \DUMP_0/dump_state_0/timer_start_RNO  (.A(
        \DUMP_0/dump_state_0/N_88 ), .B(\DUMP_0/dump_state_0/cs4 ), .Y(
        \DUMP_0/dump_state_0/timer_start_RNO_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_98  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_150_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_95_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_98_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_118  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_61_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_39_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_118_Y ));
    DFN1E1 \scalestate_0/OPENTIME[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[14]_net_1 ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i22_mux ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[13]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m38 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[18]  (.A(
        \top_code_0_dds_configdata[1] ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_502 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[18] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_107  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_15_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_112_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_107_Y ));
    AX1C \scalestate_0/necount_inc_0/XOR2_5_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount_inc_0/inc_5_net ), .C(
        \scalestate_0/necount[6]_net_1 ), .Y(
        \scalestate_0/necount1[6] ));
    MX2 \PLUSE_0/bri_timer_0/count[7]/U0  (.A(\PLUSE_0/count_2[7] ), 
        .B(\PLUSE_0/bri_timer_0/count_n7 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[7]/Y ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_16  (.A(
        \timer_top_0/dataout[11] ), .B(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_16_Y ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/ADD_20x20_slow_I19_Y_5 )
        );
    NOR2B \top_code_0/relay_on_RNO[5]  (.A(\top_code_0/N_814 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[5]_net_1 ));
    AND3 \scalestate_0/necount_inc_0/fAND2_8_inst  (.A(
        \scalestate_0/necount_inc_0/incb_2_net ), .B(
        \scalestate_0/necount_inc_0/inc_5_net ), .C(
        \scalestate_0/necount_inc_0/inc_10_net ), .Y(
        \scalestate_0/necount_inc_0/Rcout_9_net ));
    DFN1E1 \scalestate_0/CUTTIME90[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[11]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[3]  (.D(
        \DUMP_0/dump_coder_0/para4_4[3]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[3]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_19  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ), .C(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .Y(
        \timer_top_0/timer_0/N_16 ));
    AO1 \PLUSE_0/bri_state_0/cs_RNIVNCA1[14]  (.A(
        \PLUSE_0/bri_state_0/N_142 ), .B(
        \PLUSE_0/bri_state_0/cs[10]_net_1 ), .C(
        \PLUSE_0/bri_state_0/cs[14]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/N_144 ));
    NOR2 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        );
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[3]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[5] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_10_0  (.A(\xd_in[4] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout_0[4] ));
    DFN1 \DUMP_OFF_1/off_on_timer_0/count[2]  (.D(
        \DUMP_OFF_1/off_on_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/count_4[2] ));
    NOR3C \DUMP_OFF_0/off_on_coder_0/i_RNO[1]  (.A(
        \DUMP_OFF_0/off_on_coder_0/i_0_2[1] ), .B(
        \DUMP_OFF_0/off_on_coder_0/i_0_1[1] ), .C(
        bri_dump_sw_0_reset_out), .Y(
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[1] ));
    DFN1E1 \plusestate_0/PLUSETIME[4]  (.D(\top_code_0_plusedata[4] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[4]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_41_i ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[7]_net_1 ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_13  (.A(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .B(
        \timer_top_0/dataout[11] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_13_Y ));
    DFN1 \top_code_0/scan_start_ret_3  (.D(\top_code_0/N_108 ), .CLK(
        GLA_net_1), .Q(\top_code_0/N_108_reto ));
    DFN1E1 \top_code_0/pd_pluse_data[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[14] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[13]  (.D(
        \top_code_0_state_1ms_data[13] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[13]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[10]  (.A(
        \DDS_0/dds_state_0/para[10]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_290 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[10] ));
    DFN0C0 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[3] ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add )
        , .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[3] ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[0]  (.D(
        \DUMP_0/dump_coder_0/para4_4[0]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[0]_net_1 ));
    NOR3B \top_code_0/noise_start_ret_2_RNO  (.A(
        \top_code_0/un1_xa_10_2 ), .B(\top_code_0/N_332 ), .C(
        \top_code_0/N_165 ), .Y(\top_code_0/un1_xa_13 ));
    AO1 \scalestate_0/timecount_ret_90_RNO  (.A(
        \scalestate_0/CUTTIME180[8]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[8] ), .Y(
        \scalestate_0/timecount_20_iv_2[8] ));
    AX1C \CAL_0/cal_div_0/un3_count_I_12  (.A(
        \CAL_0/cal_div_0/count[3]_net_1 ), .B(
        \CAL_0/cal_div_0/DWACT_FINC_E[0] ), .C(
        \CAL_0/cal_div_0/count[4]_net_1 ), .Y(\CAL_0/cal_div_0/I_12 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m44 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[15] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[13]  (.D(
        \top_code_0_pd_pluse_data[13] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[13]_net_1 ));
    NOR2A \noisestate_0/timecount_1_RNO[15]  (.A(\noisestate_0/N_72 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[15] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_RNO[0]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[0] ));
    OA1B \syn_md_module_1/syn_md_0/count_RNO[2]  (.A(
        \syn_md_module_1/syn_md_0/N_25 ), .B(
        \syn_md_module_1/syn_md_0/count_n2_i_0 ), .C(
        \syn_md_module_1/syn_md_0/N_50 ), .Y(
        \syn_md_module_1/syn_md_0/count_RNO[2]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[8] ));
    DFN1E1 \top_code_0/state_1ms_lc[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/state_1ms_lc_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_lc[2] ));
    NOR2B \state_1ms_0/timecount_RNO_1[17]  (.A(
        \state_1ms_0/CUTTIME[17]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/timecount_8[17] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIPTS7[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[0]_net_1 ), .B(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_0[0] ));
    AO1A \scalestate_0/timecount_ret_41_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[2]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[2] ), .Y(
        \scalestate_0/timecount_20_iv_0[2] ));
    NOR2B \scalestate_0/timecount_ret_35_RNO_0  (.A(
        \scalestate_0/CUTTIMEI90[9]_net_1 ), .B(\scalestate_0/N_252 ), 
        .Y(\scalestate_0/CUTTIMEI90_m[9] ));
    NOR3C \scalestate_0/timecount_ret_5_RNO_1  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[2]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[2] ));
    NOR2B \topctrlchange_0/interupt_RNO  (.A(\topctrlchange_0/N_8 ), 
        .B(net_27), .Y(\topctrlchange_0/interupt_RNO_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[10] ));
    DFN1 \timer_top_0/timer_0/timedata[2]  (.D(
        \timer_top_0/timer_0/timedata_4[2] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[2]_net_1 ));
    OR2 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_8  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_8_net_1 )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI2909[4]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_22[0] ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_38  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[3]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[5] ));
    MX2A \scalestate_0/M_pulse_RNO_0  (.A(\scalestate_0/M_pulse8_NE ), 
        .B(\scalestate_0/M_pulse_net_1 ), .S(\scalestate_0/N_1181 ), 
        .Y(\scalestate_0/N_745 ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIPTG52[5]  (.A(
        \DUMP_0/dump_timer_0/count_c4 ), .B(\DUMP_0/count_0[5] ), .Y(
        \DUMP_0/dump_timer_0/count_c5 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[18]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_53 ), .Y(
        \timer_top_0/timer_0/timedata_4[18] ));
    NOR3C \scalestate_0/timecount_ret_1_RNO_6  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[5]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[5] ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_AGB  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_0_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_2_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_1_Y ), .Y(
        \timer_top_0/timer_0/cmp_result ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIJQII[5]  (.A(
        \DUMP_0/dump_coder_0/para4[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_5[0] ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNI7ACG[0]  (.A(
        \DUMP_0/dump_coder_0/para2[0]_net_1 ), .B(\DUMP_0/count_1[0] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_0_0[0] ));
    AO1A \scalestate_0/timecount_ret_41_RNO_2  (.A(
        \scalestate_0/N_1069 ), .B(\scalestate_0/CUTTIME90[2]_net_1 ), 
        .C(\scalestate_0/CUTTIMEI90_m[2] ), .Y(
        \scalestate_0/timecount_20_iv_4[2] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[9] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[20]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[20]_net_1 ));
    NOR2A \scalestate_0/strippluse_RNO_1[11]  (.A(\scalestate_0/N_431 )
        , .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[11] ));
    DFN1E1 \plusestate_0/PLUSETIME[5]  (.D(\top_code_0_plusedata[5] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[5]_net_1 ));
    DFN1 \state_1ms_0/timecount[1]  (.D(
        \state_1ms_0/timecount_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[1] ));
    OR3 \scalestate_0/timecount_ret_91_RNO  (.A(
        \scalestate_0/PLUSETIME90_m[8] ), .B(
        \scalestate_0/DUMPTIME_m[8] ), .C(
        \scalestate_0/S_DUMPTIME_m[8] ), .Y(
        \scalestate_0/timecount_20_iv_6[8] ));
    DFN1 \scalestate_0/strippluse[2]  (.D(
        \scalestate_0/strippluse_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[2] ));
    IOIN_IB \ADC_pad[3]/U0/U1  (.YIN(\ADC_pad[3]/U0/NET1 ), .Y(
        \ADC_c[3] ));
    DFN1E1 \top_code_0/scaleddsdiv[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[3] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[4]  (.A(
        \scalestate_0_strippluse[4] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[4] ));
    IOIN_IB \xa_pad[15]/U0/U1  (.YIN(\xa_pad[15]/U0/NET1 ), .Y(
        \xa_c[15] ));
    MX2 \nsctrl_choice_0/dumponoff_rst_RNO_0  (.A(net_33_0), .B(
        top_code_0_noise_rst_0), .S(top_code_0_n_s_ctrl_0), .Y(
        \nsctrl_choice_0/dumponoff_rst_5 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[1]  (
        .D(\s_acq_change_0_s_acqnum[1] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[1]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m48  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_47 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_48 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_49 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg_RNID0TG[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[2]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_2 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_56_i ));
    NOR3C \DDS_0/dds_timer_0/count_0_sqmuxa  (.A(dds_change_0_dds_conf)
        , .B(\DDS_0/dds_state_0_state_over ), .C(dds_change_0_dds_rst), 
        .Y(\DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[5]  (.A(
        \state_1ms_0_timecount[5] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_217 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[9] ));
    AND2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_26  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_44_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[2] )
        );
    DFN1E0 \DUMP_0/dump_coder_0/para4[11]  (.D(
        \DUMP_0/dump_coder_0/para4_4[11]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[11]_net_1 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[4]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[4] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[4]_net_1 ));
    OR2A \scalestate_0/dump_start_RNO_1  (.A(\scalestate_0/N_1196 ), 
        .B(\scalestate_0/N_1241 ), .Y(\scalestate_0/N_1167 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m43_3 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_2_RNO_1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[3]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3_0 )
        );
    DFN1E1 \plusestate_0/PLUSETIME[7]  (.D(\top_code_0_plusedata[7] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[7]_net_1 ));
    XA1 \DUMP_0/off_on_timer_1/count_RNO[1]  (.A(\DUMP_0/count_0[1] ), 
        .B(\DUMP_0/count_0[0] ), .C(
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_1/count_n1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[10]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNISL1G[4]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[4]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_4[0] ));
    NOR2A \scalestate_0/timecount_20_iv_4_RNO_0[4]  (.A(
        \scalestate_0/CUTTIME90[4]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[4] ));
    DFN1E1 \noisestate_0/dectime[13]  (.D(\top_code_0_noisedata[13] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[13]_net_1 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[11]  (.A(\s_acq_change_0/N_81 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[11]_net_1 ));
    OR2A \scalestate_0/CS_i_RNI7I7A[0]  (.A(
        \scalestate_0/CS_i[0]_net_1 ), .B(\scalestate_0/CS[16]_net_1 ), 
        .Y(\scalestate_0/N_1212 ));
    AX1C \PLUSE_0/bri_timer_0/count_RNO[7]  (.A(\PLUSE_0/count_2[6] ), 
        .B(\PLUSE_0/bri_timer_0/count_c5 ), .C(\PLUSE_0/count_2[7] ), 
        .Y(\PLUSE_0/bri_timer_0/count_n7 ));
    MX2B \noisestate_0/timecount_1_RNO[11]  (.A(\noisestate_0/N_68 ), 
        .B(\noisestate_0/N_193 ), .S(\noisestate_0/N_228 ), .Y(
        \noisestate_0/timecount_5[11] ));
    NOR2B \noisestate_0/n_acq_RNO  (.A(\noisestate_0/N_129 ), .B(
        top_code_0_noise_rst), .Y(\noisestate_0/n_acq_RNO_net_1 ));
    NOR3C \ClockManagement_0/clk_div500_0/count_RNIKKD24[0]  (.A(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_5 ), .B(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_4 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_6 ), .Y(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ));
    DFN1E1 \state_1ms_0/CUTTIME[17]  (.D(
        \top_code_0_state_1ms_data[1] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_380 ), .Q(\state_1ms_0/CUTTIME[17]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[4]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[4] ));
    NOR2B \scalestate_0/timecount_20_iv_4_RNO[11]  (.A(
        \scalestate_0/CUTTIMEI90[11]_net_1 ), .B(\scalestate_0/N_252 ), 
        .Y(\scalestate_0/CUTTIMEI90_m[11] ));
    OR3 OR3_0 (.A(DUMP_OFF_1_dump_off), .B(DUMP_OFF_0_dump_off), .C(
        DUMP_0_dump_off), .Y(dumpoff_c));
    MX2 \bri_dump_sw_0/pluse_start_RNO_0  (.A(plusestate_0_off_test), 
        .B(scalestate_0_pluse_start), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/pluse_start_5 ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m46_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[15]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[14] )
        , .Y(\DDS_0/dds_state_0/N_493 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[3]  (.A(
        \state_1ms_0_timecount[3] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_227 ));
    DFN1E1 \scanstate_0/dectime[5]  (.D(\top_code_0_scandata[5] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[5]_net_1 ));
    NOR2B \PLUSE_0/qq_state_0/stateover_0_sqmuxa_i_o3  (.A(
        \PLUSE_0/i_9[0] ), .B(bri_dump_sw_0_reset_out), .Y(
        \PLUSE_0/qq_state_0/cs4 ));
    MX2 \DSTimer_0/dump_sustain_timer_0/data_RNO_0[3]  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[3]_net_1 ), .B(
        \top_code_0_dump_sustain_data[3] ), .S(\DSTimer_0/AND2_0_Y ), 
        .Y(\DSTimer_0/dump_sustain_timer_0/N_27 ));
    DFN1E1 \scalestate_0/timecount_ret_64  (.D(
        \scalestate_0/timecount_20_iv_6[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[13] ));
    NOR2B \state_1ms_0/timecount_RNO[7]  (.A(\state_1ms_0/N_74 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[7]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[19]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[19]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_506 ));
    DFN1 \ClockManagement_0/clk_10k_0/count[7]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[7] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[7]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI7M6T[15]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[15]_net_1 ), .B(
        \sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_15[0] ));
    OR3 \state_1ms_0/timecount_RNO_1[15]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[15] ), .B(
        \state_1ms_0/CUTTIME_m[15] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[15] ), .Y(
        \state_1ms_0/timecount_8[15] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_43  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_43_Y ));
    DFN1 \scalestate_0/necount[3]  (.D(
        \scalestate_0/necount_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[3]_net_1 ));
    NOR3C \bridge_div_0/clk_4f_RNO_0  (.A(
        \bridge_div_0/clear1_n17_NE[0] ), .B(pd_pulse_en_c), .C(
        \bridge_div_0/un1_count_i[0] ), .Y(
        \bridge_div_0/clk_4f_1_sqmuxa ));
    IOPAD_IN \xa_pad[17]/U0/U0  (.PAD(xa[17]), .Y(\xa_pad[17]/U0/NET1 )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m46_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[13] ));
    DFN1 \DUMP_0/dump_timer_0/count[4]  (.D(
        \DUMP_0/dump_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_1[4] ));
    NOR2A \scalestate_0/timecount_ret_61_RNO_0  (.A(
        \scalestate_0/ACQTIME[12]_net_1 ), .B(\scalestate_0/N_1065 ), 
        .Y(\scalestate_0/ACQTIME_m[12] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[2]_net_1 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[7]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[16]  (.A(
        \DDS_0/dds_state_0/para[16]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_294 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[16] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIM9121[8]  (.A(
        \sd_acq_top_0/count_1[8] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[8]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_18[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_3[0] ));
    NOR3C \scalestate_0/timecount_ret_71_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[15]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[15] ));
    NOR2A \PLUSE_0/qq_timer_1/count_RNO[0]  (.A(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ), .B(
        \PLUSE_0/count_7[0] ), .Y(\PLUSE_0/qq_timer_1/count_n0 ));
    AND2A \PLUSE_0/bri_coder_0/half_0_I_9  (.A(\PLUSE_0/count_2[6] ), 
        .B(\PLUSE_0/half_para[6] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[2] ));
    DFN1 \bri_dump_sw_0/dumpoff_ctr  (.D(
        \bri_dump_sw_0/dumpoff_ctr_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_dumpoff_ctr));
    NOR2A \DDS_0/dds_state_0/para_reg_69_e_1  (.A(top_code_0_dds_load), 
        .B(top_code_0_dds_choice), .Y(\DDS_0/dds_state_0/N_538_1 ));
    DFN1E1 \scalestate_0/M_NUM[5]  (.D(\top_code_0_scaledatain[5] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[5]_net_1 ));
    DFN1 \plusestate_0/off_test  (.D(
        \plusestate_0/off_test_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        plusestate_0_off_test));
    DFN1E1 \noisestate_0/acqtime[11]  (.D(\top_code_0_noisedata[11] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[11]_net_1 ));
    IOTRI_OB_EB \pulse_start_pad/U0/U1  (.D(pulse_start_c), .E(VCC), 
        .DOUT(\pulse_start_pad/U0/NET1 ), .EOUT(
        \pulse_start_pad/U0/NET2 ));
    AO1C \plusestate_0/CS_RNO_0[8]  (.A(\plusestate_0/CS[2]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst), .Y(
        \plusestate_0/CS_srsts_i_0[8] ));
    MX2 \bridge_div_0/clk_4f/U0  (.A(\bridge_div_0/clk_4f_5 ), .B(
        \bridge_div_0/clk_4f ), .S(\bridge_div_0/clk_4f_1_sqmuxa ), .Y(
        \bridge_div_0/clk_4f/Y ));
    NOR2A \scalestate_0/timecount_ret_61_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[12]_net_1 ), .B(\scalestate_0/N_1089 )
        , .Y(\scalestate_0/S_DUMPTIME_m[12] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m56  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_55 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_56 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_57 ));
    DFN1 \DUMP_OFF_1/off_on_coder_0/i[0]  (.D(
        \DUMP_OFF_1/off_on_coder_0/i_RNO_4[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/i_4[0] ));
    DFN1 \ClockManagement_0/clk_10k_0/count[4]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[4] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[4]_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_2[8]  (.A(
        \state_1ms_0/M_DUMPTIME[8]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[8] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[8] ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_1_inst  (.A(
        \scalestate_0/necount[0]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .Y(
        \scalestate_0/necount1[1] ));
    DFN1E1 \scalestate_0/NE_NUM[10]  (.D(\top_code_0_scaledatain[10] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[10]_net_1 ));
    OR2A \scalestate_0/CS_RNIOAT91[12]  (.A(\scalestate_0/N_1069 ), .B(
        \scalestate_0/N_252 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_4 ));
    DFN1E1 \scalestate_0/DUMPTIME[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[10]_net_1 ));
    MX2 \scalestate_0/CS_RNO_0[20]  (.A(\scalestate_0/CS[20]_net_1 ), 
        .B(\scalestate_0/CS[9]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1232 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[1]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[1]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_8[1] ));
    IOPAD_IN \xa_pad[4]/U0/U0  (.PAD(xa[4]), .Y(\xa_pad[4]/U0/NET1 ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BFF1_0_inst  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[4] ));
    XOR2 \CAL_0/cal_div_0/count_RNIO0VJ[0]  (.A(
        \CAL_0/cal_div_0/count[0]_net_1 ), .B(\CAL_0/cal_para_out[0] ), 
        .Y(\CAL_0/cal_div_0/clear_n4_0 ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_1  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_1_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_3_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1D_0_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_1_Y ));
    MX2 \scanstate_0/timecount_1_RNO[6]  (.A(\scanstate_0/N_64 ), .B(
        \scanstate_0/timecount_cnst[2] ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[6] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[10]  (.A(
        \scalestate_0/ACQ180_NUM[10]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[10]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_458 ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[1]  (.D(
        \DUMP_0/dump_coder_0/para5_4[1] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[1]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m41_2 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_15[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[13]_net_1 ), 
        .B(\pd_pluse_top_0/count[13] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_13[0] ));
    AOI1 \DUMP_0/off_on_state_0/cs_RNIHHE1[1]  (.A(DUMP_0_dump_off), 
        .B(\DUMP_0/i_1[1] ), .C(\DUMP_0/off_on_state_0/cs[1]_net_1 ), 
        .Y(\DUMP_0/off_on_state_0/N_42_i ));
    NOR2B \DUMP_0/dump_timer_0/count_RNIT0UP1[4]  (.A(
        \DUMP_0/dump_timer_0/count_c3 ), .B(\DUMP_0/count_1[4] ), .Y(
        \DUMP_0/dump_timer_0/count_c4 ));
    DFN1E0 \DDS_0/dds_state_0/para[5]  (.D(\DDS_0/dds_state_0/N_81 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[5]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m41_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[18] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_60_i ));
    NOR2B \state_1ms_0/rt_sw_RNO  (.A(\state_1ms_0/N_153 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(\state_1ms_0/rt_sw_RNO_3 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m200  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_201 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m44_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_3  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_3_Y ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_7  (.A(
        \scalestate_0/M_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_7_Y ));
    OR2A \scalestate_0/CS_RNI83I81[5]  (.A(\scalestate_0/N_1210 ), .B(
        \scalestate_0/timecount_8_sqmuxa_i_0 ), .Y(
        \scalestate_0/N_1089 ));
    NOR2A \scanstate_0/timecount_1_RNO[10]  (.A(\scanstate_0/N_68 ), 
        .B(\scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[10] ));
    IOPAD_TRI \relay_on_pad[5]/U0/U0  (.D(\relay_on_pad[5]/U0/NET1 ), 
        .E(\relay_on_pad[5]/U0/NET2 ), .PAD(relay_on[5]));
    OR2A \plusestate_0/sw_acq1_RNO  (.A(top_code_0_pluse_rst), .B(
        \plusestate_0/N_120 ), .Y(\plusestate_0/sw_acq1_RNO_net_1 ));
    IOIN_IB \xwe_pad/U0/U1  (.YIN(\xwe_pad/U0/NET1 ), .Y(xwe_c));
    IOPAD_IN \ADC_pad[7]/U0/U0  (.PAD(ADC[7]), .Y(\ADC_pad[7]/U0/NET1 )
        );
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[0]  (.D(
        \top_code_0_halfdata_0[0] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[0] ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_0  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_12_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_2_Y ), .C(
        \timer_top_0/dataout[9] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_0_Y ));
    NOR2B \dds_change_0/dds_rst_RNO_3  (.A(top_code_0_pluse_rst), .B(
        \top_code_0_change[1] ), .Y(\dds_change_0/ddsrstin3_m ));
    NOR3C \scalestate_0/timecount_ret_19_RNO_0  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[8]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[8] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[10] ));
    OR3 \scalestate_0/timecount_ret_65_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[13] ), .B(
        \scalestate_0/OPENTIME_TEL_m[13] ), .C(
        \scalestate_0/timecount_20_iv_4[13] ), .Y(
        \scalestate_0/timecount_20_iv_8[13] ));
    DFN1E1 \scalestate_0/PLUSETIME180[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[8]_net_1 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_40  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[2] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_30  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_103_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_91_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_30_Y ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[18]  (.D(
        \top_code_0_dds_configdata[1] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[18]_net_1 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[4]  (.A(
        \timer_top_0/state_switch_0/N_220 ), .B(
        \timer_top_0/state_switch_0/N_221 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[4] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[4]_net_1 ));
    DFN1P0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]  (
        .D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_e0 ), 
        .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .PRE(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        );
    NOR3A \PLUSE_0/bri_state_0/cs_RNO_0[5]  (.A(
        \PLUSE_0/bri_state_0/cs[4]_net_1 ), .B(\PLUSE_0/i_3[2] ), .C(
        \PLUSE_0/i_8[1] ), .Y(\PLUSE_0/bri_state_0/csse_4_0_a4_0_0 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m229  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_228 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_229 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_230 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m103  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_102 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_103 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_104 ));
    AO1A \scalestate_0/timecount_ret_29_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[1]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[1] ), .Y(
        \scalestate_0/timecount_20_iv_0[1] ));
    DFN1 \state_1ms_0/timecount[14]  (.D(
        \state_1ms_0/timecount_RNO[14]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[14] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_110  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_110_Y ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[9]  (.D(
        \DUMP_0/dump_coder_0/para4_4[9]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[9]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNO_net_1 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_net_1 ));
    MX2 \s_acq_change_0/s_load_5  (.A(top_code_0_s_load), .B(
        scalestate_0_load_out), .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_load_5_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[11]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[11] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[11] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[10]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[10] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m89  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_86 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_89 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_90 ));
    DFN1E1 \scalestate_0/timecount_ret_75  (.D(
        \scalestate_0/timecount_20_iv_8[5]_net_1 ), .CLK(GLA_net_1), 
        .E(\scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[5] ));
    NOR2B \scalestate_0/necount_RNO[10]  (.A(\scalestate_0/N_740 ), .B(
        top_code_0_scale_rst_3), .Y(
        \scalestate_0/necount_RNO[10]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIOQP6[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[0]_net_1 ), .B(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_0[0] ));
    OR3 \top_code_0/cal_load_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/N_204 ));
    DFN1 \top_code_0/scale_start_ret_3  (.D(\top_code_0/N_110 ), .CLK(
        GLA_net_1), .Q(\top_code_0/N_110_reto ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_11_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_14_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net )
        , .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_11_net ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[3]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[3] ));
    MX2 \top_code_0/scan_start_ret_2_RNILFTL  (.A(
        \top_code_0/top_code_0_scan_start_reto ), .B(
        \top_code_0/un1_xa_10_reto ), .S(\top_code_0/N_108_reto ), .Y(
        \top_code_0/N_796_reto ));
    INV \syn_md_module_1/syn_md_edge_detect_0/sig_r1_RNO  (.A(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_net_1 ), .Y(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_i ));
    NOR2A \state_1ms_0/timecount_RNO_5[5]  (.A(
        \state_1ms_0/CS[5]_net_1 ), .B(
        \state_1ms_0/PLUSETIME[5]_net_1 ), .Y(
        \state_1ms_0/PLUSETIME_i_m[5] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_56  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_56_Y ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[2]  (.A(
        \s_acq_change_0/s_acqnum_5[2] ), .B(
        \s_acq_change_0_s_acqnum[2] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_72 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[12]  (.A(
        \ClockManagement_0/long_timer_0/count_c11 ), .B(
        \ClockManagement_0/long_timer_0/count[12]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n12 ));
    NOR3B \top_code_0/k2_RNO_2  (.A(\top_code_0/N_13 ), .B(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_1 ), .C(
        \top_code_0/N_154 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_3_net_1 ));
    OA1C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[10]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 ), .B(
        \pd_pluse_top_0/i_1[3] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_179 ));
    XA1 \DUMP_OFF_0/off_on_timer_0/count_RNO[1]  (.A(
        \DUMP_OFF_0/count_3[1] ), .B(\DUMP_OFF_0/count_3[0] ), .C(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_n1 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_21  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[4] )
        );
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[11]  (.D(
        \top_code_0_pd_pluse_data[11] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[11]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[2]  (.D(
        \DUMP_0/dump_coder_0/para2_4[2]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[2]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[7] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_58_i ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_8  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_2_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_11_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_0_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_8_Y ));
    AO1A \scalestate_0/timecount_ret_34_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/S_DUMPTIME[9]_net_1 ), .C(
        \scalestate_0/timecount_20_iv_1[9] ), .Y(
        \scalestate_0/timecount_20_iv_6[9] ));
    DFN1 \nsctrl_choice_0/dumpoff_ctr  (.D(
        \nsctrl_choice_0/dumpoff_ctr_RNO_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_dumpoff_ctr));
    DFN1 \topctrlchange_0/interupt  (.D(
        \topctrlchange_0/interupt_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        interupt_c));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i16_mux ));
    XA1A \timer_top_0/timer_0/Timer_Cmp_0/AND2_2  (.A(
        \timer_top_0/dataout[11] ), .B(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_27_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_2_Y ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIK1DM[6]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8 ), .B(
        \s_acq_change_0_s_stripnum[6] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_6 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[13]  (.A(
        \noisestate_0_timecount[13] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_190 ));
    AO1C \state_1ms_0/CS_RNO_0[4]  (.A(\state_1ms_0/CS[3]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[4] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[1] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i16_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_153  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_153_Y ));
    DFN1E1 \scalestate_0/CUTTIMEI90[17]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[17]_net_1 )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[5] ));
    DFN1E1 \scalestate_0/ACQTIME[8]  (.D(\top_code_0_scaledatain[8] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[8]_net_1 ));
    DFN1E1 \top_code_0/n_acqnum[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[6] ));
    DFN1E1 \scanstate_0/acqtime[7]  (.D(\top_code_0_scandata[7] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[7]_net_1 ));
    NOR2B \scalestate_0/off_test_RNO  (.A(\scalestate_0/N_726 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/off_test_RNO_1_net_1 ));
    NOR2A \state_1ms_0/un1_PLUSECYCLE13_i_a2_0_0  (.A(
        \top_code_0_state_1ms_lc[2] ), .B(\top_code_0_state_1ms_lc[1] )
        , .Y(\state_1ms_0/un1_PLUSECYCLE13_i_a2_0_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[4]  (.D(
        \top_code_0_n_acqnum_2[4] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[4]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[7]_net_1 ));
    MX2 \scalestate_0/CS_RNO_0[12]  (.A(\scalestate_0/CS[12]_net_1 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1226 ));
    DFN1 \timer_top_0/timer_0/timedata[12]  (.D(
        \timer_top_0/timer_0/timedata_4[12] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_65  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_90_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_38_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_65_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_69  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_69_Y ));
    OAI1 \scanstate_0/CS_RNIDEQ01[2]  (.A(\scanstate_0/CS[4]_net_1 ), 
        .B(\scanstate_0/CS[2]_net_1 ), .C(net_33_0), .Y(
        \scanstate_0/N_233 ));
    DFN1 \top_code_0/relay_close[1]  (.D(
        \top_code_0/relay_close_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[1] ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[3]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_37_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[3] ));
    NOR2A \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk_RNO_0  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/un1_clk_wire )
        );
    NOR2B \scalestate_0/s_acqnum_1_RNO[1]  (.A(\scalestate_0/N_548 ), 
        .B(top_code_0_scale_rst_5), .Y(
        \scalestate_0/s_acqnum_1_RNO[1]_net_1 ));
    DFN1 \state_1ms_0/CS[4]  (.D(\state_1ms_0/CS_RNO_3[4] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[4]_net_1 ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_6  (.A(
        \scalestate_0/NE_NUM[7]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_7 ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m46_2 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i6_mux ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNITSPL5[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_9[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_8[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_14[0] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[2]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[2] ));
    DFN1E1 \top_code_0/noisedata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[7] ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y ));
    IOPAD_TRI \dumpon_pad/U0/U0  (.D(\dumpon_pad/U0/NET1 ), .E(
        \dumpon_pad/U0/NET2 ), .PAD(dumpon));
    DFN1E1 \state_1ms_0/PLUSETIME[0]  (.D(
        \top_code_0_state_1ms_data[0] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[0]_net_1 ));
    OR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_1  (
        .A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[1]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_0 ));
    OA1 \sd_acq_top_0/sd_sacq_state_0/en2_RNO  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_203 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/en2_0_0_o3_0 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/en2_RNO_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_3[14]  (.A(
        \state_1ms_0/CUTTIME[14]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[14] ));
    DFN1E1 \scalestate_0/S_DUMPTIME[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[1]_net_1 ));
    DFN1 \topctrlchange_0/sw_acq1  (.D(
        \topctrlchange_0/sw_acq1_RNO_1_net_1 ), .CLK(GLA_net_1), .Q(
        sw_acq1_c));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[10]  (.A(
        \timer_top_0/state_switch_0/N_250 ), .B(
        \timer_top_0/state_switch_0/N_251 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[10] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[10]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNI9CCG[1]  (.A(
        \DUMP_0/dump_coder_0/para2[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_1[0] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[11]  (.A(
        \scalestate_0_strippluse[11] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[11] ));
    DFN1E0 \DDS_0/dds_state_0/para[32]  (.D(\DDS_0/dds_state_0/N_27 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[32]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[3]  (.A(
        \plusestate_0_timecount[3] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_229 ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_33  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[0]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[0] ));
    AO1C \scanstate_0/CS_RNO_0[4]  (.A(\scanstate_0/CS[3]_net_1 ), .B(
        timer_top_0_clk_en_scan), .C(net_33_0), .Y(
        \scanstate_0/CS_srsts_i_0[4] ));
    MX2 \noisestate_0/timecount_1_RNO_0[9]  (.A(
        \noisestate_0/acqtime[9]_net_1 ), .B(
        \noisestate_0/dectime[9]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_66 ));
    NOR2B \DUMP_OFF_0/off_on_timer_0/count_RNI5MNA[1]  (.A(
        \DUMP_OFF_0/count_3[0] ), .B(\DUMP_OFF_0/count_3[1] ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_c1 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_30  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_42_i ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[6] )
        );
    DFN1E1 \scalestate_0/timecount_ret_38  (.D(
        \scalestate_0/timecount_20_iv_8[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[3] ));
    NOR2B \DUMP_ON_0/off_on_coder_0/i_RNO[0]  (.A(OR2_1_Y), .B(OR2_2_Y)
        , .Y(\DUMP_ON_0/off_on_coder_0/i_RNO_5[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m280  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_281 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[9]  (.A(
        \top_code_0_s_acqnum_2[9] ), .B(\scalestate_0_s_acqnum[9] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[9] ));
    AO1 \scalestate_0/timecount_ret_2_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[6]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[6] ), 
        .Y(\scalestate_0/timecount_20_iv_3[6] ));
    NOR3A \scalestate_0/M_pulse_RNIJJN9_0  (.A(
        \scalestate_0/CS[15]_net_1 ), .B(
        \scalestate_0/necount_LE_M_net_1 ), .C(
        \scalestate_0/M_pulse_net_1 ), .Y(
        \scalestate_0/timecount_17_sqmuxa_1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[2]  (
        .D(\s_acq_change_0_s_acqnum[2] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[2]_net_1 )
        );
    DFN1E1 \top_code_0/halfdata[4]  (.D(\GPMI_0_dataout_0[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[4] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_21  (.A(
        \timer_top_0/dataout[15] ), .B(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_21_Y ));
    NOR2B \DDS_0/dds_timer_0/count_RNIA6NG[3]  (.A(
        \DDS_0/dds_timer_0/count_c2 ), .B(\DDS_0/count[3] ), .Y(
        \DDS_0/dds_timer_0/count_c3 ));
    AO1 \timer_top_0/state_switch_0/dataout_RNO[16]  (.A(
        \state_1ms_0_timecount[16] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .C(
        \timer_top_0/state_switch_0/N_266 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[16]_net_1 ));
    NOR3B \top_code_0/n_divnum_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/N_339 ), .C(\top_code_0/N_152 ), .Y(
        \top_code_0/n_divnum_1_sqmuxa ));
    MX2 \DSTimer_0/dump_sustain_timer_0/data_RNO_0[2]  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[2]_net_1 ), .B(
        \top_code_0_dump_sustain_data[2] ), .S(\DSTimer_0/AND2_0_Y ), 
        .Y(\DSTimer_0/dump_sustain_timer_0/N_26 ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_15  (.A(\PLUSE_0/half_para[2] ), 
        .B(\PLUSE_0/count_8[2] ), .Y(\PLUSE_0/bri_coder_0/N_3 ));
    OA1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[5]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 ), .B(
        \sd_acq_top_0/i_5[2] ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs[1]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_216 ));
    MX2B \top_code_0/scale_rst_0_0_RNI66353  (.A(
        top_code_0_scale_rst_0), .B(\top_code_0/N_159 ), .S(
        \top_code_0/N_321 ), .Y(\top_code_0/N_801 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m183  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_184 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/ADD_20x20_slow_I19_Y_6 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[19] ));
    OR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIVO7HK1[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10 ));
    XA1 \ClockManagement_0/clk_div500_0/clk_5K_RNO  (.A(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .B(
        \ClockManagement_0/clk_div500_0_clk_5K ), .C(net_27), .Y(
        \ClockManagement_0/clk_div500_0/clk_5K_RNO_net_1 ));
    AND3 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_25  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[2] )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[1] )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] )
        );
    NOR2A \PLUSE_0/bri_coder_0/half_0_I_16  (.A(\PLUSE_0/count_8[0] ), 
        .B(\PLUSE_0/half_para[0] ), .Y(\PLUSE_0/bri_coder_0/N_4 ));
    NOR2B \topctrlchange_0/interupt_RNO_2  (.A(scalestate_0_tetw_pluse)
        , .B(\top_code_0_change[0] ), .Y(\topctrlchange_0/interin2_m ));
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_29  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[0] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[1] ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[2] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[3] ));
    OA1B \noisestate_0/CS_RNO[6]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[6]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[6] )
        , .Y(\noisestate_0/CS_RNO[6]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[4]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[3] ), 
        .Y(\DDS_0/dds_state_0/N_315 ));
    NOR2B \state_1ms_0/timecount_RNO_3[12]  (.A(
        \state_1ms_0/CUTTIME[12]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/CUTTIME_m[12] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[9]_net_1 ));
    AX1C \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_5_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/count_1[6] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[6] ));
    OA1C \top_code_0/sd_sacq_load_RNO  (.A(\top_code_0/N_195 ), .B(
        top_code_0_sd_sacq_load), .C(\top_code_0/N_310 ), .Y(
        \top_code_0/N_102 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[5]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[5] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_5_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[5] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_26  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_62_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_117_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_26_Y ));
    AO1 \DUMP_0/dump_state_0/cs_RNIEUTM[6]  (.A(
        \DUMP_0/dump_state_0/N_203 ), .B(
        \DUMP_0/dump_state_0_on_start ), .C(
        \DUMP_0/dump_state_0/cs[6]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_166 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i8_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_58  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_11_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_5_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_58_Y ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_58_i ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_110_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_1_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_404 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[13]  (.D(
        \top_code_0_state_1ms_data[13] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[13]_net_1 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_8  (.A(\xd_in[6] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[6] ));
    DFN1 \pd_pluse_top_0/pd_pluse_coder_0/i[1]  (.D(\i_0_0[1] ), .CLK(
        ddsclkout_c), .Q(\i_6[1] ));
    DFN1E1 \top_code_0/scaledatain[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[14] ));
    AO1A \scalestate_0/timecount_ret_38_RNO_2  (.A(
        \scalestate_0/N_1069 ), .B(\scalestate_0/CUTTIME90[3]_net_1 ), 
        .C(\scalestate_0/CUTTIMEI90_m[3] ), .Y(
        \scalestate_0/timecount_20_iv_4[3] ));
    DFN1E1 \top_code_0/scalechoice_0[0]  (.D(\GPMI_0_dataout[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0_0[0] ));
    NOR2A \scalestate_0/un1_PLUSETIME9032_i_a2_0  (.A(
        \top_code_0_scalechoice_0[2] ), .B(
        \top_code_0_scalechoice_0[3] ), .Y(\scalestate_0/N_66 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[7]  (.A(
        \scalestate_0/ACQ180_NUM[7]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[7]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_455 ));
    AO1B \scalestate_0/CS_RNIR1C72_1[18]  (.A(\scalestate_0/N_1310 ), 
        .B(timer_top_0_clk_en_scale_0), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/un1_CS6_33_1 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[14]  (.A(
        \ClockManagement_0/long_timer_0/count_c13 ), .B(
        \ClockManagement_0/long_timer_0/count[14]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n14 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[30]  (.A(
        \DDS_0/dds_state_0/N_516 ), .B(\DDS_0/dds_state_0/N_515 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[30] ), .Y(
        \DDS_0/dds_state_0/N_169 ));
    AO1B \plusestate_0/CS_RNO_0[1]  (.A(\plusestate_0/CS_i[0]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_srsts_i_0[1] ));
    NOR2B \state_1ms_0/timecount_RNO_6[10]  (.A(
        \state_1ms_0/PLUSETIME[10]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[10] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/ADD_20x20_slow_I19_Y )
        );
    NOR2B \s_acq_change_0/s_acqnum_RNO[8]  (.A(\s_acq_change_0/N_78 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[8]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i10_mux ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m43_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[16] ));
    OR3 \scalestate_0/timecount_ret_45_RNIJ1I  (.A(
        \scalestate_0/timecount_20_0_iv_0_reto[16] ), .B(
        \scalestate_0/OPENTIME_TEL_m_reto[16] ), .C(
        \scalestate_0/timecount_20_0_iv_4_reto[16] ), .Y(
        \scalestate_0_timecount[16] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/ADD_20x20_slow_I19_Y_6 )
        );
    DFN1 \plusestate_0/CS[7]  (.D(\plusestate_0/CS_RNO_0[7] ), .CLK(
        GLA_net_1), .Q(\plusestate_0/CS[7]_net_1 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[7]  (.A(\s_acq_change_0/N_63 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[7]_net_1 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[5]  (.D(\top_code_0_scaledatain[5] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[5]_net_1 ));
    NOR3A \top_code_0/scandata_1_sqmuxa_0_a2  (.A(
        \top_code_0/scandata_1_sqmuxa_0_a2_0_net_1 ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_142 ), .Y(
        \top_code_0/scandata_1_sqmuxa ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[9]_net_1 ));
    NOR2B \scalestate_0/CS_RNO[14]  (.A(\scalestate_0/N_1227 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[14]_net_1 ));
    AND3 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3_I_8  (
        .A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIKJJB2[2]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/N_2 ));
    XA1 \DDS_0/dds_timer_0/count_RNO[1]  (.A(\DDS_0/count[1] ), .B(
        \DDS_0/count[0] ), .C(\DDS_0/dds_timer_0/count_0_sqmuxa_net_1 )
        , .Y(\DDS_0/dds_timer_0/count_n1 ));
    NOR3B \bridge_div_0/count_RNIIQOM7[4]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[4]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIIQOM7[4]_net_1 ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_44  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[9] ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[10] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i20_mux ));
    NOR3A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_2[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_6[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_9[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_12[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_11[4] ));
    NOR3B \top_code_0/n_acqnum_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/n_acqnum_1_sqmuxa_0_a2_0 ), .C(\top_code_0/N_152 ), 
        .Y(\top_code_0/n_acqnum_1_sqmuxa ));
    OA1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNILKJB2[3]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNILKJB2[3]_net_1 )
        );
    NOR3C \ClockManagement_0/clk_div500_0/un1_count_1_I_43  (.A(
        \ClockManagement_0/clk_div500_0/count[2]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[3]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_1[0] ), 
        .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[5]  (.A(
        \DUMP_0/dump_timer_0/count_c4 ), .B(\DUMP_0/count_0[5] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n5 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[12]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_68_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[14]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[14] ));
    AO1C \PLUSE_0/bri_coder_0/half_0_I_22  (.A(\PLUSE_0/half_para[3] ), 
        .B(\PLUSE_0/count_8[3] ), .C(\PLUSE_0/bri_coder_0/N_5 ), .Y(
        \PLUSE_0/bri_coder_0/N_10 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[8] ));
    IOTRI_OB_EB \relay_close_pad[6]/U0/U1  (.D(\relay_close_c[6] ), .E(
        VCC), .DOUT(\relay_close_pad[6]/U0/NET1 ), .EOUT(
        \relay_close_pad[6]/U0/NET2 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[5]_net_1 ));
    NOR3B \scalestate_0/CUTTIME90_472_e  (.A(\scalestate_0/N_62 ), .B(
        \scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/N_1685 ));
    IOTRI_OB_EB \sw_acq2_pad/U0/U1  (.D(sw_acq2_c), .E(VCC), .DOUT(
        \sw_acq2_pad/U0/NET1 ), .EOUT(\sw_acq2_pad/U0/NET2 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI6U971[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_6[0] ));
    OR3 \scalestate_0/timecount_ret_48_RNIJ2I  (.A(
        \scalestate_0/timecount_20_0_iv_0_reto[17] ), .B(
        \scalestate_0/OPENTIME_TEL_m_reto[17] ), .C(
        \scalestate_0/timecount_20_0_iv_4_reto[17] ), .Y(
        \scalestate_0_timecount[17] ));
    OR2 \top_code_0/relay_close_1_sqmuxa_0_o2_1  (.A(\xa_c[3] ), .B(
        \top_code_0/N_144 ), .Y(\top_code_0/N_154 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m224  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_225 ));
    DFN1 \top_code_0/relay_on[2]  (.D(
        \top_code_0/relay_on_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[2] ));
    NOR2A \scalestate_0/timecount_ret_68_RNO_4  (.A(
        \scalestate_0/CUTTIME90[14]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[14] ));
    NOR2A \pd_pluse_top_0/pd_pluse_state_0/cs_RNI6H1P[1]  (.A(
        \pd_pluse_top_0/i_1[2] ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[1]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_187 ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIMRFH[7]  (.A(
        \DUMP_0/dump_coder_0/para3[7]_net_1 ), .B(\DUMP_0/count_0[7] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_7[0] ));
    XOR2 \bridge_div_0/count_5_I_14  (.A(\bridge_div_0/N_2 ), .B(
        \bridge_div_0/count_RNIJROM7[5]_net_1 ), .Y(
        \bridge_div_0/count_5[5] ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_18[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_17[10] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_19[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_21[10] ));
    DFN1 \scalestate_0/dump_sustain_ctrl  (.D(
        \scalestate_0/dump_sustain_ctrl_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(scalestate_0_dump_sustain_ctrl));
    DFN1 \top_code_0/relay_close[3]  (.D(
        \top_code_0/relay_close_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[3] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[15]  (.A(
        \plusestate_0_timecount[15] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_189 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m272  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_273 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m77  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_76 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_77 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_78 ));
    DFN1 \top_code_0/relay_on[1]  (.D(
        \top_code_0/relay_on_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[1] ));
    INV \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[0]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/un1_noise_addr_0_i[0] )
        );
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI8EBK[5]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9 ), .B(
        \s_acq_change_0_s_stripnum[5] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_5 ));
    DFN1E1 \scalestate_0/CUTTIME90[16]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[16]_net_1 ));
    DFN1 \state_1ms_0/timecount[10]  (.D(
        \state_1ms_0/timecount_RNO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[10] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[10]_net_1 ));
    NOR2B \dds_change_0/dds_rst_RNO  (.A(\dds_change_0/N_5 ), .B(
        net_27), .Y(\dds_change_0/dds_rst_RNO_net_1 ));
    XO1 \scalestate_0/M_pulse_RNO_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/M_NUM[8]_net_1 ), .C(\scalestate_0/M_pulse8_7 ), 
        .Y(\scalestate_0/M_pulse8_NE_3 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[1]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[1] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[1]_net_1 )
        );
    NOR2B \s_acq_change_0/s_stripnum_RNO[8]  (.A(\s_acq_change_0/N_64 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[8]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_data[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[8] ));
    AO1A \PLUSE_0/bri_state_0/cs_RNO[12]  (.A(clk_4f_en), .B(
        \PLUSE_0/bri_state_0/cs_i_0[12] ), .C(
        \PLUSE_0/bri_state_0/N_183 ), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_0[12] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_5  (.A(\ADC_c[5] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n2 ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[0]_net_1 ));
    AOI1 \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[8]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 ), .B(
        \sd_acq_top_0/i_5[2] ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs[7]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_221 ));
    DFN1E1 \scalestate_0/timecount_ret_11  (.D(
        \scalestate_0/timecount_20_iv_7[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[7] ));
    DFN1 \noisestate_0/state_over_n  (.D(
        \noisestate_0/state_over_n_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        noisestate_0_state_over_n));
    OR3 \scalestate_0/timecount_ret_25_RNIL7I  (.A(
        \scalestate_0/timecount_20_iv_3_reto[11] ), .B(
        \scalestate_0/timecount_20_iv_2_reto[11] ), .C(
        \scalestate_0/timecount_20_iv_6_reto[11] ), .Y(
        \scalestate_0/timecount_20_iv_9_reto[11] ));
    OA1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11_0 ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_10_0 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9_0 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_28  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_18_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_96_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_28_Y ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_2  (.A(\xd_in[12] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[12] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m53  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_52 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_53 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_54 ));
    OA1B \scanstate_0/CS_RNO[1]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[1]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[1] ), 
        .Y(\scanstate_0/CS_RNO_2[1] ));
    OR2B \DDS_0/dds_state_0/cs_RNIVMGF[2]  (.A(
        \DDS_0/dds_state_0/cs[2]_net_1 ), .B(\DDS_0/i[2] ), .Y(
        \DDS_0/dds_state_0/N_227 ));
    MX2 \PLUSE_0/bri_timer_0/count[4]/U0  (.A(\PLUSE_0/count_8[4] ), 
        .B(\PLUSE_0/bri_timer_0/count_n4 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[4]/Y ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_39_i ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIEEFQ1[20]  (.A(
        \sd_acq_top_0/count[20] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[20]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_19[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_1[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_158  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_80_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_166_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_158_Y ));
    DFN1E1 \state_1ms_0/PLUSETIME[2]  (.D(
        \top_code_0_state_1ms_data[2] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[2]_net_1 ));
    OA1B \plusestate_0/CS_RNO[4]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[4]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[4] )
        , .Y(\plusestate_0/CS_RNO_0[4]_net_1 ));
    DFN1E1 \top_code_0/s_addchoice_0[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_0[4] ));
    MX2 \PLUSE_0/bri_coder_0/i[0]/U0  (.A(\PLUSE_0/i_8[0] ), .B(
        pulse_start_c), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_coder_0/i[0]/Y ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIBIII[1]  (.A(
        \DUMP_0/dump_coder_0/para4[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_1[0] ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_62_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_0 ));
    DFN1E1 \noisestate_0/acqtime[14]  (.D(\top_code_0_noisedata[14] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[14]_net_1 ));
    NOR2B \scalestate_0/necount_LE_NE_RNIMS0L  (.A(
        \scalestate_0/N_1267 ), .B(top_code_0_scale_rst_3), .Y(
        \scalestate_0/timecount_11_sqmuxa ));
    NOR3B 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa_0_a2  
        (.A(\top_code_0_pd_pluse_choice[1] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/N_12 ), .C(
        \top_code_0_pd_pluse_choice[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_10  (.A(\ADC_c[0] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(\Signal_Noise_Acq_0/n_adc_1_10 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[6]_net_1 ));
    DFN1E1 \plusestate_0/PLUSETIME[1]  (.D(\top_code_0_plusedata[1] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[1]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_51_RNO_0  (.A(
        \scalestate_0/CUTTIME180[18]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[18] ));
    DFN1E1 \scalestate_0/OPENTIME[8]  (.D(\top_code_0_scaledatain[8] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[8]_net_1 ));
    NOR3B \top_code_0/s_periodnum_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/s_periodnum_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_152 ), .Y(\top_code_0/s_periodnum_1_sqmuxa ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_8  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/NE_NUM[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_8_Y ));
    NOR2B \ClockManagement_0/clk_10k_0/clk_5M_reg2_RNO  (.A(net_27), 
        .B(\ClockManagement_0/clk_10k_0/clk_5M_reg1_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/clk_5M_reg2_RNO_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_2[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_2[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_1[10] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_11[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_17[10] ));
    IOTRI_OB_EB \dumpoff_pad/U0/U1  (.D(dumpoff_c), .E(VCC), .DOUT(
        \dumpoff_pad/U0/NET1 ), .EOUT(\dumpoff_pad/U0/NET2 ));
    OR2A \topctrlchange_0/sw_acq2_RNO  (.A(net_27), .B(
        \topctrlchange_0/N_9 ), .Y(\topctrlchange_0/sw_acq2_RNO_3 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIVD6T[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_11[0] ));
    NOR2A \top_code_0/un1_xa_13_0_a2_0  (.A(\xa_c[2] ), .B(\xa_c[4] ), 
        .Y(\top_code_0/N_332 ));
    RAM512X18 #( .MEMORYFILE("RAM_R0C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R0C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_0_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_0_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_0_net ));
    NOR2 \top_code_0/scaleload_RNO_1  (.A(\top_code_0/N_174 ), .B(
        \top_code_0/N_159 ), .Y(\top_code_0/N_304 ));
    XA1A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_4[4]  (.A(
        \pd_pluse_top_0/count_6[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[0]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_0[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_8[4] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[21]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[22]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_512 ));
    NOR3B \top_code_0/state_1ms_data_1_sqmuxa_0_a2_1  (.A(
        \top_code_0/N_333 ), .B(\xa_c[4] ), .C(\xa_c[2] ), .Y(
        \top_code_0/state_1ms_data_1_sqmuxa_0_a2_1_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m99  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_100 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_37_i ));
    DFN1 \scalestate_0/necount[9]  (.D(
        \scalestate_0/necount_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[9]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m41_5 ));
    NOR3B \plusestate_0/sw_acq1_RNO_1  (.A(\plusestate_0/N_302 ), .B(
        \plusestate_0/N_301 ), .C(\plusestate_0/CS[8]_net_1 ), .Y(
        \plusestate_0/N_298 ));
    NOR2A \top_code_0/scandata_1_sqmuxa_0_a2_0  (.A(net_27), .B(
        \top_code_0/N_157 ), .Y(
        \top_code_0/scandata_1_sqmuxa_0_a2_0_net_1 ));
    OR3 \PLUSE_0/qq_coder_0/i_reg10_NE_3[0]  (.A(
        \PLUSE_0/qq_coder_0/i_reg10_2[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_0/i_reg10_3[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_0/i_reg10_NE_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_NE_3[0]_net_1 ));
    DFN1E1 \state_1ms_0/PLUSETIME[1]  (.D(
        \top_code_0_state_1ms_data[1] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[1]_net_1 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_2_RNO_0  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3_0 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I2_un1_CO1 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_3 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[3] ));
    NOR2B \DDS_0/dds_timer_0/count_RNIF2TK[4]  (.A(
        \DDS_0/dds_timer_0/count_c3 ), .B(\DDS_0/count[4] ), .Y(
        \DDS_0/dds_timer_0/count_c4 ));
    DFN1 \timer_top_0/state_switch_0/dataout[11]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[11]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[11] ));
    DFN1C0 \PLUSE_0/bri_coder_0/i[0]/U1  (.D(
        \PLUSE_0/bri_coder_0/i[0]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/i_8[0] ));
    DFN1 \noisestate_0/sw_acq2  (.D(\noisestate_0/sw_acq2_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(noisestate_0_sw_acq2));
    NOR2B \top_code_0/state_1ms_start_ret_1_RNI05H21  (.A(
        \top_code_0/N_797_reto ), .B(\top_code_0/net_27_reto ), .Y(
        top_code_0_scale_start));
    NOR2A \GPMI_0/tri_state_0/dataout_1_12_0  (.A(\xd_in[2] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout_0[2] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[9]_net_1 ));
    AND2 \ClockManagement_0/clk_div500_0/un1_count_1_I_53  (.A(
        \ClockManagement_0/clk_div500_0/count[4]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_1_1[0] )
        );
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[12]  (.A(
        \plusestate_0_timecount[12] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_259 ));
    DFN1E1 \plusestate_0/PLUSETIME[3]  (.D(\top_code_0_plusedata[3] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[3]_net_1 ));
    NOR3A \scalestate_0/necount_cmp_1/NOR3A_0  (.A(
        \scalestate_0/necount_cmp_1/OR2A_0_Y ), .B(
        \scalestate_0/necount_cmp_1/AO1C_2_Y ), .C(
        \scalestate_0/NE_NUM[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/NOR3A_0_Y ));
    AX1C \timer_top_0/timer_0/un2_timedata_I_26  (.A(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[4] ), .C(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .Y(
        \timer_top_0/timer_0/I_26_0 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m41_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[18] ));
    OR3 \scalestate_0/timecount_ret_63_RNIJ7I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[13] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[13] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[13] ), .Y(
        \scalestate_0_timecount[13] ));
    DFN1E1 \noisestate_0/dectime[3]  (.D(\top_code_0_noisedata[3] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[3]_net_1 ));
    DFN1 \bri_dump_sw_0/phase_ctr  (.D(
        \bri_dump_sw_0/phase_ctr_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_phase_ctr));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI0ICH[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_11[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_4_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_5_net ), 
        .B(\pd_pluse_top_0/count_1[5] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[5] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[9]  (.A(\DDS_0/dds_state_0/N_289 )
        , .B(\DDS_0/dds_state_0/N_288 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[9] ), .Y(
        \DDS_0/dds_state_0/N_14 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI6Q301[9]  (
        .A(\pd_pluse_top_0/count_0[9] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[9]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_6[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_5[0] ));
    IOPAD_TRI \relay_on_pad[8]/U0/U0  (.D(\relay_on_pad[8]/U0/NET1 ), 
        .E(\relay_on_pad[8]/U0/NET2 ), .PAD(relay_on[8]));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[2]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \top_code_0_dds_configdata[1] ), .Y(\DDS_0/dds_state_0/N_485 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[5]  (.A(\s_acq_change_0/N_75 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[5]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_1[0]_net_1 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_0[0]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_2[0]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]_net_1 ));
    DFN1 \DUMP_OFF_0/off_on_state_0/cs[1]  (.D(
        \DUMP_OFF_0/off_on_state_0/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/off_on_state_0/cs[1]_net_1 ));
    MX2B \top_code_0/k1_RNO_0  (.A(k1_c), .B(\xa_c[0] ), .S(
        \top_code_0/N_11 ), .Y(\top_code_0/N_807 ));
    DFN1 \state_1ms_0/CS[3]  (.D(\state_1ms_0/CS_RNO_3[3] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[3]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i10_mux ));
    RAM512X18 #( .MEMORYFILE("RAM_R15C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R15C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_15_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_15_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_0_net )
        );
    NOR2B \DDS_0/dds_timer_0/count_RNI6BHC[2]  (.A(
        \DDS_0/dds_timer_0/count_c1 ), .B(\DDS_0/count[2] ), .Y(
        \DDS_0/dds_timer_0/count_c2 ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_21  (.A(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[3] ));
    XA1A \syn_md_module_1/syn_md_0/count_RNO_0[3]  (.A(
        \syn_md_module_1/syn_md_0/N_18 ), .B(
        \syn_md_module_1/syn_md_0/count[3]_net_1 ), .C(
        top_code_0_scale_rst_1), .Y(\syn_md_module_1/syn_md_0/N_22 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m223  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_224 ));
    AO1B \DDS_0/dds_state_0/state_over_RNO  (.A(
        \DDS_0/dds_state_0_state_over ), .B(\DDS_0/dds_state_0/N_451 ), 
        .C(\DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/state_over_RNO_net_1 ));
    DFN1 \top_code_0/scan_rst  (.D(
        \top_code_0/scan_rst_RNIMNCI3_net_1 ), .CLK(GLA_net_1), .Q(
        net_33));
    OR2 \top_code_0/cal_data_1_sqmuxa_0_o2  (.A(\top_code_0/N_149 ), 
        .B(\xa_c[0] ), .Y(\top_code_0/N_165 ));
    MX2B \plusestate_0/timecount_1_RNO[6]  (.A(\plusestate_0/N_77 ), 
        .B(\plusestate_0/N_223 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[6] ));
    NOR2A \noisestate_0/timecount_1_RNO[13]  (.A(\noisestate_0/N_70 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[13] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNINBV25[12]  (.A(
        \ClockManagement_0/long_timer_0/count_c11 ), .B(
        \ClockManagement_0/long_timer_0/count[12]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c12 ));
    NOR2B \state_1ms_0/timecount_RNO[3]  (.A(\state_1ms_0/N_70 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[3]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIC6HP9[3]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_13[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_12[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_16[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_19[0] ));
    DFN1 \s_acq_change_0/s_stripnum[9]  (.D(
        \s_acq_change_0/s_stripnum_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[9] ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[8]  (.A(
        \s_acq_change_0/s_stripnum_5[8] ), .B(
        \s_acq_change_0_s_stripnum[8] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_64 ));
    OR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_4 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_5 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1_net_1 )
        );
    DFN1 \DUMP_OFF_1/off_on_coder_0/i[1]  (.D(
        \DUMP_OFF_1/off_on_coder_0/i_RNO_4[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/i_4[1] ));
    DFN1 \scanstate_0/CS_i_0[0]  (.D(\scanstate_0/CS_i_0_RNO_0[0] ), 
        .CLK(GLA_net_1), .Q(\scanstate_0/CS_li[0] ));
    OR3 \bridge_div_0/count_RNIVP8P3[4]  (.A(
        \bridge_div_0/un1_count_NE_0[0] ), .B(
        \bridge_div_0/un1_count_0[0] ), .C(
        \bridge_div_0/un1_count_NE_1[0] ), .Y(
        \bridge_div_0/un1_count_i[0] ));
    DFN1E1 \scalestate_0/DUMPTIME[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[12]_net_1 ));
    DFN1E1 \bridge_div_0/datahalf[2]  (.D(\top_code_0_scaleddsdiv[2] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/datahalf[2]_net_1 ));
    MX2 \top_code_0/relay_on_RNO_0[5]  (.A(\relay_on_c[5] ), .B(
        \GPMI_0_dataout[5] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_814 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[11]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[11] ));
    XA1 \DUMP_0/off_on_timer_1/count_RNO[4]  (.A(
        \DUMP_0/off_on_timer_1/count_9_0 ), .B(\DUMP_0/count_0[4] ), 
        .C(\DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_1/count_n4 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_3  (.A(
        \timer_top_0/dataout[7] ), .B(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_5_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_3_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[6] ));
    NOR2 \scalestate_0/reset_out_RNO_5  (.A(
        \scalestate_0/CS[12]_net_1 ), .B(\scalestate_0/CS[6]_net_1 ), 
        .Y(\scalestate_0/un1_CS6_39_i_a3_0 ));
    IOIN_IB \xa_pad[4]/U0/U1  (.YIN(\xa_pad[4]/U0/NET1 ), .Y(\xa_c[4] )
        );
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7_132_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ));
    MX2 \scalestate_0/CS_RNO_0[16]  (.A(\scalestate_0/CS[16]_net_1 ), 
        .B(\scalestate_0/CS[15]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1229 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[12]_net_1 ));
    AO1C \scalestate_0/necount_cmp_0/AO1C_2  (.A(
        \scalestate_0/necount[4]_net_1 ), .B(
        \scalestate_0/M_NUM[4]_net_1 ), .C(
        \scalestate_0/necount[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/AO1C_2_Y ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[4] ), .CLK(
        GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 ));
    NOR3A \DUMP_0/dump_coder_0/i_RNO_3[3]  (.A(
        \DUMP_0/dump_coder_0/i_0_0_a2_1[3] ), .B(
        \DUMP_0/dump_coder_0/un1_count_4_10[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_11[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_6[3] ));
    DFN1E1 \scalestate_0/timecount_ret_94  (.D(
        \scalestate_0/un1_timecount_2_sqmuxa_7 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/un1_timecount_2_sqmuxa_7_reto ));
    DFN1 \ClockManagement_0/clk_10k_0/count[0]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[0] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[0]_net_1 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[10]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_0[10] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[10]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[5]  (.A(
        \scanstate_0_timecount[5] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_216 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_27  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[4] )
        , .B(\s_acq_change_0_s_stripnum[8] ), .C(
        \s_acq_change_0_s_stripnum[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4 ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_8  (.A(
        \top_code_0_sigtimedata[8] ), .B(
        \ClockManagement_0/long_timer_0/count[8]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_8 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_14  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] )
        );
    NOR3C \sd_acq_top_0/sd_sacq_state_0/cs_RNO[14]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[13]_net_1 ), .B(
        \sd_acq_top_0/i[10] ), .C(\sd_acq_top_0/sd_sacq_state_0/cs4 ), 
        .Y(\sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[14] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[7]  (.A(
        \scalestate_0/s_acqnum_7[7] ), .B(\scalestate_0_s_acqnum[7] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_554 ));
    OR2A \scalestate_0/sw_acq2_RNO  (.A(top_code_0_scale_rst_3), .B(
        \scalestate_0/N_541 ), .Y(\scalestate_0/sw_acq2_RNO_1 ));
    OR2A \top_code_0/state_1ms_rst_n_0_0_RNI848T5  (.A(net_27), .B(
        \top_code_0/N_800 ), .Y(
        \top_code_0/state_1ms_rst_n_0_0_RNI848T5_net_1 ));
    DFN1E1 \top_code_0/bri_datain[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[10] ));
    AND2 \scalestate_0/necount_inc_0/AND2_8_inst  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/inc_8_net ));
    NOR3B \timer_top_0/timer_0/time_up_RNIMPL21  (.A(
        \timer_top_0/state_switch_0_state_over_n ), .B(
        \timer_top_0/state_switch_0_state_start ), .C(
        \timer_top_0/timer_0_time_up ), .Y(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ));
    AO1 \scalestate_0/timecount_RNO_2[21]  (.A(
        \scalestate_0/CUTTIMEI90[21]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[21] ), .Y(
        \scalestate_0/timecount_20_0_iv_1[21] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[14]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[13] )
        , .Y(\DDS_0/dds_state_0/N_461 ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_4  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_10_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_9_Y ), .C(
        \timer_top_0/dataout[3] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_4_Y ));
    DFN1 \syn_md_module_1/syn_md_0/count[0]  (.D(
        \syn_md_module_1/syn_md_0/count_RNO_0[0]_net_1 ), .CLK(
        GLA_net_1), .Q(\syn_md_module_1/syn_md_0/count[0]_net_1 ));
    XO1 \scalestate_0/M_pulse_RNO_8  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/M_NUM[6]_net_1 ), .C(\scalestate_0/M_pulse8_5 ), 
        .Y(\scalestate_0/M_pulse8_NE_1 ));
    OR2 \scalestate_0/CS_RNI6F271[2]  (.A(\scalestate_0/N_1203 ), .B(
        \scalestate_0/N_1197 ), .Y(\scalestate_0/un1_CS_20 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_64_i ));
    INV \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[0]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/un1_noise_addr_1_i[0] )
        );
    NOR2A \top_code_0/state_1ms_start_ret_2_RNO_0  (.A(
        \top_code_0/N_329 ), .B(\top_code_0/N_140 ), .Y(
        \top_code_0/un1_xa_4_0_a2_1 ));
    DFN1 \top_code_0/relay_on[6]  (.D(
        \top_code_0/relay_on_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[6] ));
    DFN1E1 \top_code_0/bri_datain[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[1] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[11]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[11] ));
    AOI1 \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[3]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 ), .B(
        \pd_pluse_top_0/i_1[2] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs[3]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_174 ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/count[0]  (.D(
        \DSTimer_0/dump_sustain_timer_0/count_n0 ), .CLK(clock_10khz), 
        .Q(\DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ));
    IOPAD_BI \xd_pad[10]/U0/U0  (.D(\xd_pad[10]/U0/NET1 ), .E(
        \xd_pad[10]/U0/NET2 ), .Y(\xd_pad[10]/U0/NET3 ), .PAD(xd[10]));
    OR3B \scalestate_0/CS_RNO_0[18]  (.A(\scalestate_0/N_1194 ), .B(
        timer_top_0_clk_en_scale_0), .C(
        \scalestate_0/un1_CS6_31_i_o2_0 ), .Y(\scalestate_0/N_1213 ));
    DFN1E1 \scalestate_0/PLUSETIME90[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[10]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_91  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_156_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_54_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_91_Y ));
    NOR2B \state_1ms_0/timecount_RNO_6[13]  (.A(
        \state_1ms_0/PLUSETIME[13]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[13] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_7_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_7_net ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ));
    XOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIGH7R[1]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[1]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIV7QK[12]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[12]_net_1 ), .B(
        \sd_acq_top_0/count_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_12[0] ));
    DFN1E1 \scalestate_0/DUMPTIME[3]  (.D(\top_code_0_scaledatain[3] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[3]_net_1 ));
    DFN1E1 \plusestate_0/timecount_1[4]  (.D(
        \plusestate_0/timecount_5[4] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[4] ));
    MX2 \top_code_0/relay_on_RNO_0[1]  (.A(\relay_on_c[1] ), .B(
        \GPMI_0_dataout[1] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_810 ));
    MX2 \top_code_0/relay_close_RNO_0[8]  (.A(\relay_close_c[8] ), .B(
        \GPMI_0_dataout[8] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_827 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m55  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[0] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_56 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_112  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_112_Y ));
    DFN1E1 \top_code_0/plusedata[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[10] ));
    IOPAD_TRI \calcuinter_pad/U0/U0  (.D(\calcuinter_pad/U0/NET1 ), .E(
        \calcuinter_pad/U0/NET2 ), .PAD(calcuinter));
    NOR2B \bri_dump_sw_0/off_test_RNO  (.A(\bri_dump_sw_0/off_test_5 ), 
        .B(net_27), .Y(\bri_dump_sw_0/off_test_RNO_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[23]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[24]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_301 ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI9EPB2[12]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_11 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_4 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[2]  (.D(\top_code_0_scaledatain[2] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[2]_net_1 ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_11  (.A(\PLUSE_0/count_2[7] ), 
        .B(\PLUSE_0/half_para[7] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[4] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m43 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] ));
    AO1 \scalestate_0/timecount_ret_23_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[10]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[10] ), .Y(
        \scalestate_0/timecount_20_iv_4[10] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m209  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[9] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_210 ));
    NOR3A \PLUSE_0/qq_state_0/cs_RNO[2]  (.A(\PLUSE_0/qq_state_0/cs4 ), 
        .B(\PLUSE_0/qq_state_0/N_89 ), .C(\PLUSE_0/qq_state_0/N_88 ), 
        .Y(\PLUSE_0/qq_state_0/cs_RNO_1[2]_net_1 ));
    AND2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_16[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_11[0] ));
    DFN1 \scalestate_0/necount[4]  (.D(
        \scalestate_0/necount_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[4]_net_1 ));
    NOR3A \top_code_0/dds_configdata_1_sqmuxa_0_a2  (.A(
        \top_code_0/dds_configdata_1_sqmuxa_1 ), .B(\top_code_0/N_142 )
        , .C(\top_code_0/N_155 ), .Y(
        \top_code_0/dds_configdata_1_sqmuxa ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[2]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[2] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_10[2] ));
    DFN1E1 \top_code_0/state_1ms_data[9]  (.D(\GPMI_0_dataout[9] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[9] ));
    DFN1E1 \top_code_0/sigtimedata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[6] ));
    OA1C \top_code_0/nstatechoice_RNO  (.A(\top_code_0/N_210 ), .B(
        top_code_0_nstatechoice), .C(\top_code_0/N_286 ), .Y(
        \top_code_0/N_78 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[2]  (.A(
        \scalestate_0_timecount[2] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_233 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m45_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[15]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m45_3 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_6  
        (.A(\s_acq_change_0_s_stripnum[1] ), .B(
        \s_acq_change_0_s_stripnum[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_12 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[12]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[12] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_0[12] ));
    NOR3B \PLUSE_0/bri_state_0/cs_RNIVBIV[0]  (.A(
        \PLUSE_0/bri_state_0/cs[0]_net_1 ), .B(\PLUSE_0/i_1[4] ), .C(
        \PLUSE_0/i_3[3] ), .Y(\PLUSE_0/bri_state_0/N_179 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m242  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_243 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[9] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_54_i ));
    DFN1 \scalestate_0/CS[16]  (.D(\scalestate_0/CS_RNO[16]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[16]_net_1 ));
    OA1C \top_code_0/n_s_ctrl_0_RNIURA26  (.A(\top_code_0/N_198 ), .B(
        top_code_0_n_s_ctrl_0), .C(\top_code_0/N_284 ), .Y(
        \top_code_0/N_76 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m74  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_71 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_74 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_75 ));
    AO1 \scalestate_0/timecount_ret_5_RNO_2  (.A(
        \scalestate_0/CUTTIME180[2]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[2] ), .Y(
        \scalestate_0/timecount_20_iv_2[2] ));
    DFN1 \state_1ms_0/timecount[0]  (.D(
        \state_1ms_0/timecount_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[6]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[5] ), 
        .Y(\DDS_0/dds_state_0/N_274 ));
    DFN1E1 \top_code_0/sd_sacq_choice[0]  (.D(\GPMI_0_dataout[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_choice_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_choice[0] ));
    DFN1E1 \scalestate_0/PLUSETIME180[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[9]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_27  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[4] ), .B(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .Y(
        \timer_top_0/timer_0/N_13 ));
    DFN1 \bri_dump_sw_0/tetw_pluse  (.D(
        \bri_dump_sw_0/tetw_pluse_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_tetw_pluse));
    NOR3 \DDS_0/dds_state_0/para_RNO[29]  (.A(
        \DDS_0/dds_state_0/N_484 ), .B(\DDS_0/dds_state_0/N_483 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[29] ), .Y(
        \DDS_0/dds_state_0/N_131 ));
    NOR2A \DUMP_0/off_on_timer_1/count_RNO[0]  (.A(
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ), .B(
        \DUMP_0/count_0[0] ), .Y(\DUMP_0/off_on_timer_1/count_n0 ));
    NOR3C \top_code_0/k2_RNO_1  (.A(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_3_net_1 ), .B(
        \top_code_0/un1_state_1ms_rst_n117_2_i_a2_2 ), .C(
        \top_code_0/N_11_3 ), .Y(\top_code_0/N_12 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m47  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[0] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_48 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m43_4 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[15]  (.A(
        \DDS_0/dds_state_0/para[15]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_493 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[15] ));
    OA1 \scanstate_0/CS_i_0_RNO[0]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS_li[0] ), .C(net_33_0), .Y(
        \scanstate_0/CS_i_0_RNO_0[0] ));
    MX2 \plusestate_0/timecount_1_RNO_0[11]  (.A(
        \plusestate_0/PLUSETIME[11]_net_1 ), .B(
        \plusestate_0/DUMPTIME[11]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_82 ));
    DFN1E1 \plusestate_0/PLUSETIME[6]  (.D(\top_code_0_plusedata[6] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[6]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_68_i ));
    XOR2 \DSTimer_0/dump_sustain_timer_0/start_RNO_2  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[0]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/un1_data_0 ));
    DFN1E1 \scalestate_0/timecount_ret_0  (.D(
        \scalestate_0/timecount_cnst_m_0[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_cnst_m_0_reto[6] ));
    AND3B \scalestate_0/CS_RNI270V1[4]  (.A(\scalestate_0/N_1210 ), .B(
        \scalestate_0/un1_CS_20 ), .C(\scalestate_0/N_1263 ), .Y(
        \scalestate_0/N_1241 ));
    OA1 \plusestate_0/CS_i_RNO[0]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS_i[0]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_i_RNO[0]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[19]  (.A(
        \top_code_0_dds_configdata[2] ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_506 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[19] ));
    DFN1E1 \scalestate_0/timecount_ret_54  (.D(
        \scalestate_0/timecount_20_0_iv_0[19] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_0_reto[19] ));
    NOR2B \scalestate_0/timecount_ret_8_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[3]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[3] ));
    AND3 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_1_12_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_5_net )
        , .C(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_150  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_150_Y ));
    OR3 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIOSMH2[0]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_3 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_4 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_0 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_2 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[2] ));
    DFN1E1 \scalestate_0/PLUSETIME180[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[2]_net_1 ));
    OR2B \dds_change_0/un1_change_2  (.A(\top_code_0_change[1] ), .B(
        \top_code_0_change[0] ), .Y(\dds_change_0.un1_change_2 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[2]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[2] ));
    AO1 \sd_acq_top_0/sd_sacq_state_0/cs_RNI1SAS[6]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[6]_net_1 ), .B(
        \sd_acq_top_0/i_2[4] ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_235 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_203 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIG0KE2[7]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_11[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_13[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_13[0] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_27  (.A(
        \timer_top_0/dataout[10] ), .B(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_27_Y ));
    NOR2A \timer_top_0/state_switch_0/state_start5_0_0_a2_1_0  (.A(
        top_code_0_scan_start), .B(top_code_0_noise_start), .Y(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_1_0_net_1 ));
    OR3 \scalestate_0/timecount_ret_66_RNO  (.A(
        \scalestate_0/CUTTIME180_m[14] ), .B(
        \scalestate_0/OPENTIME_m[14] ), .C(
        \scalestate_0/timecount_20_iv_3[14] ), .Y(
        \scalestate_0/timecount_20_iv_7[14] ));
    OR2A \top_code_0/dumpdata_1_sqmuxa_0_o2  (.A(\xa_c[1] ), .B(
        \xa_c[0] ), .Y(\top_code_0/N_159 ));
    AO1C \state_1ms_0/CS_RNO_0[7]  (.A(\state_1ms_0/CS[6]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[7] ));
    AND3 \scalestate_0/necount_cmp_0/AND3_1  (.A(
        \scalestate_0/necount_cmp_0/XNOR2_8_Y ), .B(
        \scalestate_0/necount_cmp_0/XNOR2_5_Y ), .C(
        \scalestate_0/necount_cmp_0/XNOR2_3_Y ), .Y(
        \scalestate_0/necount_cmp_0/AND3_1_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[9] ));
    NOR3C \scalestate_0/timecount_ret_91_RNO_0  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[8]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[8] ));
    MX2 \state1ms_choice_0/dump_start_RNO_0  (.A(
        bri_dump_sw_0_dump_start), .B(state_1ms_0_dump_start), .S(
        top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/dump_start_5 ));
    OR3 \scalestate_0/timecount_ret_11_RNIA4I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[7] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[7] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[7] ), .Y(
        \scalestate_0/timecount_20_iv_10_reto[7] ));
    DFN1E1 \top_code_0/s_addchoice_1[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_1[4] ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[4]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_12_2 ), .Y(
        \timer_top_0/timer_0/timedata_4[4] ));
    DFN1E1 \scanstate_0/acqtime[3]  (.D(\top_code_0_scandata[3] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[3]_net_1 ));
    AND2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/FND2_8_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net ), 
        .B(\pd_pluse_top_0/count_0[9] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_12_net ));
    DFN1 \bri_dump_sw_0/dump_start  (.D(
        \bri_dump_sw_0/dump_start_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_dump_start));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/TAND2_15_inst  (
        .A(\sd_acq_top_0/count_0[12] ), .B(\sd_acq_top_0/count_0[13] ), 
        .C(\sd_acq_top_0/count_0[14] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net ));
    NOR2B \state_1ms_0/timecount_RNO[4]  (.A(\state_1ms_0/N_71 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[4]_net_1 ));
    NOR2 \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[6]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/en2 ), .B(
        \pd_pluse_top_0/i_1[2] ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_185 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_11  (.A(
        \timer_top_0/dataout[16] ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_11_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_125  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_125_Y ));
    AND2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_28  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[2] ));
    NOR2A \scalestate_0/timecount_ret_91_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[8]_net_1 ), .B(\scalestate_0/N_1089 ), 
        .Y(\scalestate_0/S_DUMPTIME_m[8] ));
    NOR2A \scalestate_0/timecount_ret_23_RNO_4  (.A(
        \scalestate_0/CUTTIME90[10]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[10] ));
    DFN1E1 \scanstate_0/dectime[6]  (.D(\top_code_0_scandata[6] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[6]_net_1 ));
    MX2B \scalestate_0/soft_d_RNO_0  (.A(scalestate_0_soft_d), .B(
        \scalestate_0/N_1241 ), .S(\scalestate_0/N_1259 ), .Y(
        \scalestate_0/N_543 ));
    DFN1 \scanstate_0/sw_acq2  (.D(\scanstate_0/sw_acq2_RNO_2 ), .CLK(
        GLA_net_1), .Q(scanstate_0_sw_acq2));
    XA1 \PLUSE_0/qq_timer_0/count_RNO[1]  (.A(\PLUSE_0/count_9[1] ), 
        .B(\PLUSE_0/count_9[0] ), .C(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_0/count_n1 ));
    MX2B \plusestate_0/timecount_1_RNO[1]  (.A(\plusestate_0/N_72 ), 
        .B(\plusestate_0/N_245 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[1] ));
    AO1 \scalestate_0/timecount_ret_66_RNO_2  (.A(
        \scalestate_0/CUTTIME180_TEL[14]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[14] )
        , .Y(\scalestate_0/timecount_20_iv_3[14] ));
    NOR2B \DUMP_OFF_1/off_on_coder_0/i_RNO[0]  (.A(
        nsctrl_choice_0_dumpoff_ctr), .B(nsctrl_choice_0_dumponoff_rst)
        , .Y(\DUMP_OFF_1/off_on_coder_0/i_RNO_4[0] ));
    OR2A \DUMP_0/dump_state_0/cs_RNIEVCA[4]  (.A(
        \DUMP_0/dump_state_0/cs[4]_net_1 ), .B(\DUMP_0/i_0[3] ), .Y(
        \DUMP_0/dump_state_0/N_173 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[1]  (.D(
        \DUMP_0/dump_coder_0/para4_4[1]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[1]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[1]  (.A(
        \state_1ms_0/PLUSETIME[1]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[1] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_52_i ));
    DFN1 \scanstate_0/state_over_n  (.D(
        \scanstate_0/state_over_n_RNO_1 ), .CLK(GLA_net_1), .Q(
        scanstate_0_state_over_n));
    DFN1E1 \DDS_0/dds_state_0/para_reg[1]  (.D(
        \top_code_0_dds_configdata[0] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[1]_net_1 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[4]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[4] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_10[4] ));
    NOR3C \DUMP_0/off_on_state_0/cs_RNO[0]  (.A(
        state1ms_choice_0_reset_out), .B(\DUMP_0/i_1[0] ), .C(
        \DUMP_0/off_on_state_0/N_42_i ), .Y(
        \DUMP_0/off_on_state_0/N_36_i ));
    NOR2A \plusestate_0/timecount_1_RNO[11]  (.A(\plusestate_0/N_82 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[11] ));
    NOR2 \top_code_0/s_periodnum_1_sqmuxa_0_a2_0  (.A(
        \top_code_0/N_159 ), .B(\top_code_0/N_150 ), .Y(
        \top_code_0/s_periodnum_1_sqmuxa_0_a2_0_net_1 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[14]  (.A(
        \timer_top_0/state_switch_0/N_260 ), .B(
        \timer_top_0/state_switch_0/N_261 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[14] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[14]_net_1 ));
    DFN1E1 \plusestate_0/timecount_1[5]  (.D(
        \plusestate_0/timecount_5[5] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[5] ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[15]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[15] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[15] ));
    NOR3B \top_code_0/sd_sacq_choice_1_sqmuxa_0_a2  (.A(
        \top_code_0/N_331 ), .B(\top_code_0/N_329 ), .C(
        \top_code_0/N_163 ), .Y(\top_code_0/sd_sacq_choice_1_sqmuxa ));
    NOR2B \scalestate_0/reset_out_RNO  (.A(\scalestate_0/N_540 ), .B(
        top_code_0_scale_rst), .Y(\scalestate_0/reset_out_RNO_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m289  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_288 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_289 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_290 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/YAND2_21_inst  (
        .A(\sd_acq_top_0/count_0[15] ), .B(\sd_acq_top_0/count[16] ), 
        .C(\sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_27_net ));
    DFN1E1 \scalestate_0/S_DUMPTIME[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[5]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m304  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_303 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_304 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_305 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[11] ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_30  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[4] ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_37_i ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_15_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_20_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_14_net ));
    DFN1E1 \scalestate_0/timecount_ret_85  (.D(
        \scalestate_0/timecount_20_iv_6[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[11] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_38_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_39_i ));
    AND3 \scalestate_0/necount_cmp_0/AND3_2  (.A(
        \scalestate_0/necount_cmp_0/XNOR2_0_Y ), .B(
        \scalestate_0/necount_cmp_0/XNOR2_9_Y ), .C(
        \scalestate_0/necount_cmp_0/XNOR2_7_Y ), .Y(
        \scalestate_0/necount_cmp_0/AND3_2_Y ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[10]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[10] ));
    AO1C \PLUSE_0/bri_coder_0/half_0_I_18  (.A(\PLUSE_0/count_8[1] ), 
        .B(\PLUSE_0/half_para[1] ), .C(\PLUSE_0/bri_coder_0/N_4 ), .Y(
        \PLUSE_0/bri_coder_0/N_6 ));
    DFN1 \s_acq_change_0/s_acqnum[9]  (.D(
        \s_acq_change_0/s_acqnum_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[9] ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_6  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_24_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_12_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_9_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_6_Y ));
    NOR3C \scalestate_0/CUTTIME180_TEL_510_e  (.A(\scalestate_0/N_61 ), 
        .B(\scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 ), .C(
        \top_code_0_scalechoice_0[0] ), .Y(\scalestate_0/N_1723 ));
    DFN1 \PLUSE_0/qq_state_1/cs[1]  (.D(
        \PLUSE_0/qq_state_1/cs_RNO_2[1] ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_1/cs[1]_net_1 ));
    IOIN_IB \xa_pad[17]/U0/U1  (.YIN(\xa_pad[17]/U0/NET1 ), .Y(
        \xa_c[17] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m70  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m70_1 ));
    DFN1 \DDS_0/dds_state_0/cs[3]  (.D(
        \DDS_0/dds_state_0/cs_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n3 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3]/Y ));
    DFN1E1 \scalestate_0/CUTTIMEI90[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[8]_net_1 ));
    NOR2B \state1ms_choice_0/dump_start_RNO  (.A(
        \state1ms_choice_0/dump_start_5 ), .B(net_27), .Y(
        \state1ms_choice_0/dump_start_RNO_1 ));
    NOR3 \scalestate_0/timecount_ret_93_RNO  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_6_0 ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_6_1 ), .C(
        \scalestate_0/un1_timecount_2_sqmuxa_4 ), .Y(
        \scalestate_0/timecount_m3_e_2 ));
    NOR2A \DDS_0/dds_state_0/w_clk_reg_RNIEMPL  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/w_clk_reg_net_1 ), .Y(
        \DDS_0/dds_state_0/para_1_sqmuxa_1_0 ));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/en1_RNO  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_184 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/en1_0_i_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/en1_RNO_net_1 ));
    DFN1E1 \top_code_0/bri_datain[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[8] ));
    MX2B \scanstate_0/rt_sw_RNO_0  (.A(scanstate_0_rt_sw), .B(
        \scanstate_0/CS[5]_net_1 ), .S(\scanstate_0/N_253 ), .Y(
        \scanstate_0/N_111 ));
    DFN1E1 \top_code_0/s_addchoice_3[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_3[0] ));
    AO1 \state_1ms_0/timecount_RNO_4[7]  (.A(
        \state_1ms_0/S_DUMPTIME[7]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[7] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[7] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m43_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[16] ));
    DFN1E1 \scalestate_0/PLUSETIME90[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[8]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNIKTLJ[5]  (.A(
        \DUMP_0/dump_coder_0/para5[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_5[0] ));
    NOR3C \PLUSE_0/bri_timer_0/count_RNIVCH9[4]  (.A(
        \PLUSE_0/count_8[3] ), .B(\PLUSE_0/bri_timer_0/count_c2 ), .C(
        \PLUSE_0/count_8[4] ), .Y(\PLUSE_0/bri_timer_0/count_c4 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[2]  (.A(
        \timer_top_0/state_switch_0/N_230 ), .B(
        \timer_top_0/state_switch_0/N_231 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[2] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[2]_net_1 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[1]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[1] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_6[1] ));
    AX1C \timer_top_0/timer_0/un2_timedata_I_7  (.A(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[2]_net_1 ), .Y(
        \timer_top_0/timer_0/I_7_2 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m111  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_108 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_111 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_112 ));
    OR2A \scalestate_0/sw_acq1_RNO  (.A(top_code_0_scale_rst_3), .B(
        \scalestate_0/N_542 ), .Y(\scalestate_0/sw_acq1_RNO_0_net_1 ));
    NOR3B \top_code_0/noisedata_1_sqmuxa_0_a2  (.A(\xa_c[2] ), .B(
        \top_code_0/noisedata_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_151 ), .Y(\top_code_0/noisedata_1_sqmuxa ));
    DFN1E1 \scalestate_0/PLUSETIME180[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[4]_net_1 ));
    NOR2B \syn_md_module_1/syn_md_edge_detect_0/sig_r1_RNI92I1  (.A(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r1_i_0 ), .B(
        \syn_md_module_1/syn_md_edge_detect_0/sig_r0_net_1 ), .Y(
        \syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en ));
    XOR3 \bridge_div_0/dataall_1_I_12  (.A(\top_code_0_scaleddsdiv[1] )
        , .B(\top_code_0_scaleddsdiv[4] ), .C(
        \bridge_div_0/DWACT_ADD_CI_0_TMP[0] ), .Y(
        \bridge_div_0/dataall_1[1] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[9]  (.D(
        \top_code_0_pd_pluse_data[9] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[9]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[30]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[30]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_515 ));
    NOR2B \top_code_0/sigtimedata_1_sqmuxa_0_a2_1  (.A(
        \top_code_0/N_329 ), .B(net_27), .Y(
        \top_code_0/sigtimedata_1_sqmuxa_1 ));
    IOPAD_IN \ADC_pad[10]/U0/U0  (.PAD(ADC[10]), .Y(
        \ADC_pad[10]/U0/NET1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI4MK91[15]  (.A(
        \sd_acq_top_0/count_0[15] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[15]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_12[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_4[0] ));
    OA1A \DDS_0/dds_state_0/fq_ud_reg_RNO  (.A(
        \DDS_0/dds_state_0/N_226 ), .B(\DDS_0/dds_state_0/cs[3]_net_1 )
        , .C(\DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/fq_ud_reg_RNO_net_1 ));
    DFN1 \plusestate_0/tetw_pluse  (.D(\plusestate_0/tetw_pluse_RNO_0 )
        , .CLK(GLA_net_1), .Q(plusestate_0_tetw_pluse));
    IOTRI_OB_EB \cal_out_pad/U0/U1  (.D(cal_out_c), .E(VCC), .DOUT(
        \cal_out_pad/U0/NET1 ), .EOUT(\cal_out_pad/U0/NET2 ));
    NOR2A \scalestate_0/timecount_ret_88_RNO_1  (.A(
        \scalestate_0/DUMPTIME[10]_net_1 ), .B(\scalestate_0/N_1093 ), 
        .Y(\scalestate_0/DUMPTIME_m[10] ));
    NOR3A \scalestate_0/reset_out_RNO_4  (.A(
        \scalestate_0/un1_CS6_39_i_a3_0 ), .B(
        \scalestate_0/CS_0[11]_net_1 ), .C(\scalestate_0/CS[13]_net_1 )
        , .Y(\scalestate_0/un1_CS6_39_i_a3_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[22]  (.A(
        \top_code_0_dds_configdata[5] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_459 ), .Y(
        \DDS_0/dds_state_0/para_9_i_0_1[22] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[7] ));
    DFN1E1 \top_code_0/pluse_noise_ctrl  (.D(\top_code_0/N_86 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pluse_noise_ctrl));
    NOR3 \timer_top_0/state_switch_0/state_over_n_RNO  (.A(
        \timer_top_0/state_switch_0/N_278 ), .B(
        \timer_top_0/state_switch_0/N_279 ), .C(
        \timer_top_0/state_switch_0/state_over_n_0_i_0 ), .Y(
        \timer_top_0/state_switch_0/N_78 ));
    DFN1E1 \top_code_0/scaleddsdiv[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[1] ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[12]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_35_1 ), .Y(
        \timer_top_0/timer_0/timedata_4[12] ));
    DFN1E1 \scalestate_0/timecount_ret_45  (.D(
        \scalestate_0/timecount_20_0_iv_0[16] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_0_reto[16] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[4]  (.D(
        \top_code_0_pd_pluse_data[4] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[4]_net_1 ));
    DFN1E0C0 \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_4 ), .CLK(
        ddsclkout_c), .CLR(s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_1_sqmuxa )
        , .Q(\Signal_Noise_Acq_0/signal_acq_0/clkout ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI38T7[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_5[0] ));
    DFN1E1 \scalestate_0/CUTTIME180[17]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1661 ), .Q(\scalestate_0/CUTTIME180[17]_net_1 )
        );
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_11 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_12 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_3 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_9 )
        );
    NOR3B \noisestate_0/CS_i_0_RNIGJKN[0]  (.A(\noisestate_0/CS_li[0] )
        , .B(top_code_0_noise_rst), .C(\noisestate_0/CS[5]_net_1 ), .Y(
        \noisestate_0/timecount_cnst[4] ));
    MX2 \top_code_0/relay_on_RNO_0[8]  (.A(\relay_on_c[8] ), .B(
        \GPMI_0_dataout[8] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_817 ));
    DFN1 \DUMP_0/dump_timer_0/count[6]  (.D(
        \DUMP_0/dump_timer_0/count_n6 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[6] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m204  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_197 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_204 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[10] ));
    DFN1 \PLUSE_0/qq_state_1/cs[4]  (.D(
        \PLUSE_0/qq_state_1/cs_RNO_3[4] ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_1/cs[4]_net_1 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[6]  (.A(
        \scalestate_0_strippluse[6] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[6] ));
    DFN1 \DDS_0/dds_coder_0/i[0]  (.D(
        \DDS_0/dds_coder_0/i_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/i[0] ));
    NOR2A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[12]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_195 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_0_Y ));
    XO1 \PLUSE_0/qq_coder_0/i_reg10_NE_2[0]  (.A(\PLUSE_0/count_9[1] ), 
        .B(\PLUSE_0/qq_para3[1] ), .C(
        \PLUSE_0/qq_coder_0/i_reg10_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_NE_2[0]_net_1 ));
    DFN1 \state_1ms_0/dump_start  (.D(
        \state_1ms_0/dump_start_RNO_2_net_1 ), .CLK(GLA_net_1), .Q(
        state_1ms_0_dump_start));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_73  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_67_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_151_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_73_Y ));
    NOR3A \DUMP_0/dump_coder_0/i_RNO_2[3]  (.A(
        \DUMP_0/dump_coder_0/i_0_0_a2_3[3] ), .B(
        \DUMP_0/dump_coder_0/un1_count_4_3[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_2[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_7[3] ));
    NOR2A \PLUSE_0/qq_state_1/cs_RNO[4]  (.A(\PLUSE_0/qq_state_1/cs4 ), 
        .B(\PLUSE_0/qq_state_1/N_84 ), .Y(
        \PLUSE_0/qq_state_1/cs_RNO_3[4] ));
    NOR2A \PLUSE_0/qq_coder_1/i_RNO[3]  (.A(bri_dump_sw_0_reset_out), 
        .B(\PLUSE_0/qq_coder_1/i_reg10_NE[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/i_RNO_3[3] ));
    DFN1 \bri_dump_sw_0/pluse_start  (.D(
        \bri_dump_sw_0/pluse_start_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        pulse_start_c));
    DFN1 \timer_top_0/state_switch_0/dataout[7]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[7]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[7] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[8]  (.A(
        \scalestate_0_strippluse[8] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[8] ));
    DFN1 \s_acq_change_0/s_acqnum[10]  (.D(
        \s_acq_change_0/s_acqnum_RNO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[10] ));
    NOR2A \syn_md_module_1/syn_md_0/un1_syn_md_out_en_1_i_i_a2  (.A(
        top_code_0_scale_rst_3), .B(
        \syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en ), .Y(
        \syn_md_module_1/syn_md_0/N_52 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[14]  (.A(
        \noisestate_0_timecount[14] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_260 ));
    DFN1 \DUMP_ON_0/off_on_state_0/cs[0]  (.D(
        \DUMP_ON_0/off_on_state_0/N_36_i ), .CLK(GLA_net_1), .Q(
        DUMP_ON_0_dump_on));
    DFN1 \DDS_0/dds_coder_0/i[2]  (.D(
        \DDS_0/dds_coder_0/i_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/i[2] ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[13]  (.D(
        \top_code_0_state_1ms_data[13] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[13]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[3]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[8]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[8] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 ));
    NOR2A \DUMP_ON_0/off_on_timer_0/count_RNO[0]  (.A(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_ON_0/count_5[0] ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_n0 ));
    MX2 \scanstate_0/timecount_1_RNO_0[12]  (.A(
        \scanstate_0/acqtime[12]_net_1 ), .B(
        \scanstate_0/dectime[12]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_70 ));
    DFN1 \scalestate_0/necount[10]  (.D(
        \scalestate_0/necount_RNO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[10]_net_1 ));
    DFN1E1 \top_code_0/state_1ms_lc[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/state_1ms_lc_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_lc[0] ));
    DFN1E1 \top_code_0/pluse_lc  (.D(\top_code_0/N_84 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pluse_lc));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[4]  (.A(
        \scanstate_0_timecount[4] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_221 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO_0[15]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c12 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c14 ));
    DFN1 \scalestate_0/necount[5]  (.D(
        \scalestate_0/necount_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[5]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_62_i ));
    NOR2B \noisestate_0/soft_d_RNO  (.A(\noisestate_0/N_109 ), .B(
        top_code_0_noise_rst), .Y(\noisestate_0/soft_d_RNO_net_1 ));
    MX2 \dds_change_0/dds_rst_RNO_0  (.A(dds_change_0_dds_rst), .B(
        \dds_change_0/dds_rst_6 ), .S(\dds_change_0.un1_change_2 ), .Y(
        \dds_change_0/N_5 ));
    DFN1E1 \top_code_0/s_periodnum[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_periodnum_1_sqmuxa ), .Q(
        \top_code_0_s_periodnum[2] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[3]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[3] ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_20  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7 ), .B(
        \s_acq_change_0_s_stripnum[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_20 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[3]  (.A(
        \scalestate_0/s_acqnum_7[3] ), .B(\scalestate_0_s_acqnum[3] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_550 ));
    OR3 \state_1ms_0/timecount_RNO_1[5]  (.A(
        \state_1ms_0/timecount_8_iv_1[5] ), .B(
        \state_1ms_0/timecount_8_iv_0[5] ), .C(
        \state_1ms_0/timecount_8_iv_2[5] ), .Y(
        \state_1ms_0/timecount_8_iv[5] ));
    AO1C \scalestate_0/necount_cmp_1/AO1C_1  (.A(
        \scalestate_0/necount[7]_net_1 ), .B(
        \scalestate_0/NE_NUM[7]_net_1 ), .C(
        \scalestate_0/necount[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/AO1C_1_Y ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[6]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[6] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_6_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[6] ));
    NOR2A \scalestate_0/timecount_ret_RNIEH21  (.A(
        \scalestate_0/timecount_cnst_reto[5] ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .Y(
        \scalestate_0/timecount_cnst_m_reto[5] ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_13[3]  (.A(
        \DUMP_0/dump_coder_0/para1[9]_net_1 ), .B(\DUMP_0/count[9] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_9[0] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[15]  (.A(
        \DDS_0/dds_state_0/N_496 ), .B(\DDS_0/dds_state_0/N_495 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[15] ), .Y(
        \DDS_0/dds_state_0/N_159 ));
    MX2A \state_1ms_0/timecount_RNO_0[6]  (.A(
        \state_1ms_0/timecount_8_iv[6] ), .B(
        \state_1ms_0_timecount[6] ), .S(\state_1ms_0/CS[9]_net_1 ), .Y(
        \state_1ms_0/N_73 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[2]_net_1 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_60  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_56_i ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9_0 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[4]  (.A(\scalestate_0/N_452 ), 
        .B(\scalestate_0/ACQECHO_NUM[4]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[4] ));
    DFN1E0 \DDS_0/dds_state_0/para[35]  (.D(
        \DDS_0/dds_state_0/para_9[35] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[35]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[4]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[4] ));
    OR3 \scalestate_0/timecount_20_iv_8[11]  (.A(
        \scalestate_0/timecount_20_iv_0[11] ), .B(
        \scalestate_0/OPENTIME_TEL_m[11] ), .C(
        \scalestate_0/timecount_20_iv_4[11]_net_1 ), .Y(
        \scalestate_0/timecount_20_iv_8[11]_net_1 ));
    AO1A \scalestate_0/CS_RNIE2Q31[7]  (.A(\scalestate_0/CS[7]_net_1 ), 
        .B(top_code_0_inv_turn), .C(scalestate_0_ne_le), .Y(
        \scalestate_0/un1_CS6_31_i_o2_0 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m44  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[0] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_45 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m270  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_269 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_270 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_271 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIU7QF[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_4[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_3[0] ));
    NOR3C \ClockManagement_0/long_timer_0/timeup_RNO_0  (.A(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_12 ), .B(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_11 ), .C(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_13 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa ));
    IOPAD_BI \xd_pad[5]/U0/U0  (.D(\xd_pad[5]/U0/NET1 ), .E(
        \xd_pad[5]/U0/NET2 ), .Y(\xd_pad[5]/U0/NET3 ), .PAD(xd[5]));
    DFN1E1 \top_code_0/dds_configdata[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[11] ));
    OR3 \state_1ms_0/timecount_RNO_1[1]  (.A(
        \state_1ms_0/timecount_8_iv_1[1] ), .B(
        \state_1ms_0/timecount_8_iv_0[1] ), .C(
        \state_1ms_0/timecount_8_iv_2[1] ), .Y(
        \state_1ms_0/timecount_8[1] ));
    OR2A \scalestate_0/necount_cmp_1/OR2A_1  (.A(
        \scalestate_0/NE_NUM[2]_net_1 ), .B(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OR2A_1_Y ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_50  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_48_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[8] )
        );
    DFN1E1 \state_1ms_0/S_DUMPTIME[14]  (.D(
        \top_code_0_state_1ms_data[14] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[14]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m42_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[17] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[12]_net_1 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[6]_net_1 ));
    MX2 \scalestate_0/CS_RNO_0[7]  (.A(\scalestate_0/CS[7]_net_1 ), .B(
        \scalestate_0/CS[6]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1222 ));
    DFN1E0 \DDS_0/dds_state_0/para[31]  (.D(\DDS_0/dds_state_0/N_171 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[31]_net_1 ));
    NOR3B \PLUSE_0/qq_state_0/Q1Q8_Q2Q7_RNO  (.A(
        \PLUSE_0/qq_state_0/N_79 ), .B(\PLUSE_0/qq_state_0/cs4 ), .C(
        \PLUSE_0/qq_state_0/cs[4]_net_1 ), .Y(
        \PLUSE_0/qq_state_0/Q1Q8_Q2Q7_RNO_net_1 ));
    NOR3A \top_code_0/cal_data_1_sqmuxa_0_a2  (.A(
        \top_code_0/cal_data_1_sqmuxa_1 ), .B(\xa_c[2] ), .C(
        \top_code_0/N_155 ), .Y(\top_code_0/cal_data_1_sqmuxa ));
    IOTRI_OB_EB \relay_close_pad[0]/U0/U1  (.D(\relay_close_c[0] ), .E(
        VCC), .DOUT(\relay_close_pad[0]/U0/NET1 ), .EOUT(
        \relay_close_pad[0]/U0/NET2 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[9] ));
    DFN1E1 \scalestate_0/ACQ180_NUM[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[1]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m173  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_166 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_173 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_174 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m47_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[12] ));
    NOR2B \scalestate_0/strippluse_RNO[10]  (.A(\scalestate_0/N_569 ), 
        .B(top_code_0_scale_rst_3), .Y(
        \scalestate_0/strippluse_RNO[10]_net_1 ));
    AX1C \DUMP_0/dump_timer_0/count_RNO[11]  (.A(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_0/count[11] ), .C(\DUMP_0/dump_timer_0/N_52 ), .Y(
        \DUMP_0/dump_timer_0/count_n11 ));
    NOR2A \scanstate_0/timecount_1_RNO[13]  (.A(\scanstate_0/N_71 ), 
        .B(\scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[13] ));
    DFN1E1 \scanstate_0/dectime[9]  (.D(\top_code_0_scandata[9] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[9]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[18]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[18]_net_1 ));
    OR3 \state_1ms_0/timecount_RNO_1[10]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[10] ), .B(
        \state_1ms_0/CUTTIME_m[10] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[10] ), .Y(
        \state_1ms_0/timecount_8[10] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i8_mux ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i18_mux ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[7]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_36_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[7] ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/en2  (.D(
        \sd_acq_top_0/sd_sacq_state_0/en2_RNO_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/sd_sacq_state_0/en2_net_1 ));
    XOR2 \ClockManagement_0/clk_div500_0/un1_count_1_I_31  (.A(
        \ClockManagement_0/clk_div500_0/count[4]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] ), 
        .Y(\ClockManagement_0/clk_div500_0/I_31 ));
    IOPAD_BI \xd_pad[0]/U0/U0  (.D(\xd_pad[0]/U0/NET1 ), .E(
        \xd_pad[0]/U0/NET2 ), .Y(\xd_pad[0]/U0/NET3 ), .PAD(xd[0]));
    OA1C \top_code_0/dds_load_RNO  (.A(\top_code_0/N_200 ), .B(
        top_code_0_dds_load), .C(\top_code_0/N_276 ), .Y(
        \top_code_0/N_68 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[17]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[17]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_8_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_8_net ));
    DFN1E1 \scalestate_0/timecount_ret_65  (.D(
        \scalestate_0/timecount_20_iv_8[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[13] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[2]  (.D(
        \top_code_0_n_acqnum_2[2] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[2]_net_1 ));
    DFN1 \DUMP_OFF_1/off_on_timer_0/count[0]  (.D(
        \DUMP_OFF_1/off_on_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/count_4[0] ));
    NOR2B \scalestate_0/ACQ90_NUM_1_sqmuxa_0_a2_1  (.A(
        \top_code_0_scalechoice_0[3] ), .B(
        \top_code_0_scalechoice_0[2] ), .Y(\scalestate_0/N_67 ));
    DFN1E1 \top_code_0/state_1ms_data[7]  (.D(\GPMI_0_dataout[7] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[7] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[4]  (.D(
        \top_code_0_dds_configdata[3] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[4]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_49  (.A(
        \timer_top_0/timer_0/N_6 ), .B(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .Y(
        \timer_top_0/timer_0/I_49 ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[7]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[7] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_0[7] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m119  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_116 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_119 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_120 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m41_6 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[4]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[4] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_6[4] ));
    IOPAD_TRI \sw_acq2_pad/U0/U0  (.D(\sw_acq2_pad/U0/NET1 ), .E(
        \sw_acq2_pad/U0/NET2 ), .PAD(sw_acq2));
    NOR2B \DUMP_0/dump_state_0/cs_RNIBSCA[2]  (.A(
        \DUMP_0/dump_state_0/cs[2]_net_1 ), .B(\DUMP_0/i_0[2] ), .Y(
        \DUMP_0/dump_state_0/N_196 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m284  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_285 ));
    NOR2B \PLUSE_0/bri_state_0/en  (.A(\PLUSE_0/i_8[0] ), .B(
        bri_dump_sw_0_reset_out), .Y(\PLUSE_0/bri_state_0/en_net_1 ));
    NOR2 \top_code_0/n_acqnum_1_sqmuxa_0_a2_0_0  (.A(
        \top_code_0/N_157 ), .B(\top_code_0/N_154 ), .Y(
        \top_code_0/n_acqnum_1_sqmuxa_0_a2_0 ));
    XA1 \DSTimer_0/dump_sustain_timer_0/count_RNO[2]  (.A(
        \DSTimer_0/dump_sustain_timer_0/count_c1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[2]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_n2 ));
    NOR3B \top_code_0/un1_state_1ms_rst_n117_43_i_a2_0  (.A(\xa_c[6] ), 
        .B(\top_code_0/un1_state_1ms_rst_n117_43_i_a2_0_0_net_1 ), .C(
        \top_code_0/N_137 ), .Y(\top_code_0/N_325 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m10  
        (.A(\s_acq_change_0_s_stripnum[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[3]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i6_mux ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_23  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[5]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[1] )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIBK3A[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[8]_net_1 ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_8[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_51  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_83_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_33_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_51_Y ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNILA8D[10]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[10]_net_1 )
        , .B(\pd_pluse_top_0/count_0[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_10[0] ));
    DFN1 \DUMP_0/off_on_timer_1/count[4]  (.D(
        \DUMP_0/off_on_timer_1/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[4] ));
    NOR2B \pd_pluse_top_0/pd_pluse_coder_0/i_RNO[0]  (.A(pulse_start_c)
        , .B(net_27), .Y(\pd_pluse_top_0/pd_pluse_coder_0/i_RNO_6[0] ));
    DFN1E1 \top_code_0/scaledatain[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[9] ));
    DFN1E1 \scalestate_0/CUTTIME180[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[1]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[8]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[8] ));
    NOR2B \state1ms_choice_0/bri_cycle_RNO  (.A(
        \state1ms_choice_0/bri_cycle_5 ), .B(net_27), .Y(
        \state1ms_choice_0/bri_cycle_RNO_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m203  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_200 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_203 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_204 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_10[3]  (.A(
        \DUMP_0/dump_coder_0/para1[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_11[0] ));
    DFN1E1 \top_code_0/bri_datain[14]  (.D(\GPMI_0_dataout[14] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[14] ));
    DFN1E1 \top_code_0/s_acqnum[15]  (.D(\GPMI_0_dataout[15] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[15] ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_37_i ));
    DFN1 \noisestate_0/CS[5]  (.D(\noisestate_0/CS_RNO[5]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[5]_net_1 ));
    MX2 \topctrlchange_0/rt_sw_RNO_0  (.A(rt_sw_net_0), .B(
        \topctrlchange_0/rt_sw_6 ), .S(\dds_change_0.un1_change_2 ), 
        .Y(\topctrlchange_0/N_12 ));
    NOR2B \scalestate_0/timecount_ret_84_RNO_0  (.A(
        \scalestate_0/CUTTIME180[11]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[11] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[21]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[21]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_9_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_9_net ));
    XO1 \PLUSE_0/qq_coder_0/un1_qq_para2_NE_0[0]  (.A(
        \PLUSE_0/count_9[4] ), .B(\PLUSE_0/qq_para2[4] ), .C(
        \PLUSE_0/qq_para2[5] ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_0[0]_net_1 ));
    OA1B \state_1ms_0/CS_RNO[9]  (.A(\state_1ms_0/CS[9]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(\state_1ms_0/CS_srsts_i_0[9] ), 
        .Y(\state_1ms_0/CS_RNO_1[9] ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNIA09M3[7]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c6 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c8 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[0]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[0] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_10[0] ));
    DFN1E1 \scanstate_0/dectime[2]  (.D(\top_code_0_scandata[2] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[2]_net_1 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[14]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[14] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count[14] ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNIQ3MJ[8]  (.A(
        \DUMP_0/dump_coder_0/para5[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_8[0] ));
    DFN1E1 \top_code_0/scaleload  (.D(\top_code_0/N_96 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_scaleload));
    NOR2B \PLUSE_0/qq_state_1/stateover_0_sqmuxa_i_o3  (.A(
        \PLUSE_0/i_7[0] ), .B(bri_dump_sw_0_reset_out), .Y(
        \PLUSE_0/qq_state_1/cs4 ));
    DFN1P0 \PLUSE_0/bri_state_0/cs[12]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_0[12] ), .CLK(ddsclkout_c), .PRE(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs_i_0[12] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_4  (.A(\xd_in[10] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[10] ));
    NOR3B \scalestate_0/timecount_ret_27_RNIN9I  (.A(
        \scalestate_0/timecount_m3_e_1_reto ), .B(
        \scalestate_0/timecount_m3_e_2_reto ), .C(
        \scalestate_0/un1_timecount_2_sqmuxa_7_reto ), .Y(
        \scalestate_0/timecount_11_sqmuxa_m_reto ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[8]  (.A(
        \s_acq_change_0/s_acqnum_5[8] ), .B(
        \s_acq_change_0_s_acqnum[8] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_78 ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_1  (.A(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .B(
        \timer_top_0/dataout[1] ), .C(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_1_Y ));
    NOR3C \PLUSE_0/bri_state_0/cs_RNO_2[3]  (.A(
        \PLUSE_0/bri_state_0/cs_i_0[7] ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[13] ), .C(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_1 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_6 ));
    DFN1E1 \plusestate_0/PLUSETIME[12]  (.D(\top_code_0_plusedata[12] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[12]_net_1 ));
    OR3 \scalestate_0/timecount_ret_60_RNO  (.A(
        \scalestate_0/CUTTIME180_m[12] ), .B(
        \scalestate_0/OPENTIME_m[12] ), .C(
        \scalestate_0/timecount_20_iv_3[12] ), .Y(
        \scalestate_0/timecount_20_iv_7[12] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_13_0  (.A(\xd_in[1] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout_0[1] ));
    DFN1E1 \top_code_0/noisedata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[6] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_147  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_159_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_147_Y ));
    MX2 \scalestate_0/s_acq180_RNO_0  (.A(\scalestate_0/CS[9]_net_1 ), 
        .B(s_acq180_c), .S(\scalestate_0/un1_CS6 ), .Y(
        \scalestate_0/N_742 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[6]  (.A(
        \top_code_0_dumpdata_0[6] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[6] ));
    DFN1 \state_1ms_0/CS[5]  (.D(\state_1ms_0/CS_RNO_3[5] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[5]_net_1 ));
    DFN1E1 \top_code_0/dumpdata[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[2] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[2]  (.A(
        \DDS_0/dds_state_0/para[2]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_485 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[2] ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_15[3]  (.A(
        \DUMP_0/dump_coder_0/para1[1]_net_1 ), .B(\DUMP_0/count_1[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_1[0] ));
    OR3 \state_1ms_0/timecount_RNO_1[8]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[8] ), .B(
        \state_1ms_0/CUTTIME_m[8] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[8] ), .Y(
        \state_1ms_0/timecount_8[8] ));
    DFN1 \DUMP_0/dump_coder_0/i[7]  (.D(
        \DUMP_0/dump_coder_0/i_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i[7] ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[2]  (.A(
        \ClockManagement_0/long_timer_0/count_c1 ), .B(
        \ClockManagement_0/long_timer_0/count[2]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n2 ));
    NOR2B \scalestate_0/strippluse_RNO[1]  (.A(\scalestate_0/N_560 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[1]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m297  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_296 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_297 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_298 ));
    NOR2B \ClockManagement_0/clk_10k_0/count_RNITQ4S[5]  (.A(
        \ClockManagement_0/clk_10k_0/count[5]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[6]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_2 ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[1]  (.D(
        \top_code_0_cal_data[1] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[1] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_3  (.A(
        \timer_top_0/dataout[3] ), .B(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_3_Y ));
    IOTRI_OB_EB \relay_on_pad[5]/U0/U1  (.D(\relay_on_c[5] ), .E(VCC), 
        .DOUT(\relay_on_pad[5]/U0/NET1 ), .EOUT(
        \relay_on_pad[5]/U0/NET2 ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[0]  (.D(
        \DUMP_0/dump_coder_0/para4_4[0]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[0]_net_1 ));
    DFN1E1 \top_code_0/n_acqnum[4]  (.D(\GPMI_0_dataout_0[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[4] ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_0  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_7_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_2_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_6_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_0_Y ));
    NOR2A \scalestate_0/strippluse_RNO_1[6]  (.A(\scalestate_0/N_426 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[6] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[14]_net_1 )
        );
    NOR3A \DUMP_0/dump_coder_0/para16  (.A(\top_code_0_dump_cho_0[0] ), 
        .B(\top_code_0_dump_cho_0[2] ), .C(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para16_net_1 ));
    DFN1E1 \scalestate_0/ACQTIME[2]  (.D(\top_code_0_scaledatain_0[2] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[2]_net_1 ));
    XA1C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_11[4]  (.A(
        \pd_pluse_top_0/count[14] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[14]_net_1 ), 
        .C(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_11[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_1[4] ));
    DFN1E1 \top_code_0/acqclken  (.D(\top_code_0/N_60 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_acqclken));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_33  
        (.A(\s_acq_change_0_s_stripnum[9] ), .B(
        \s_acq_change_0_s_stripnum[10] ), .C(
        \s_acq_change_0_s_stripnum[11] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[7] )
        );
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[4]  (.A(
        \top_code_0_dumpdata_0[4] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[4] ));
    OR3 \scalestate_0/timecount_ret_61_RNO  (.A(
        \scalestate_0/ACQTIME_m[12] ), .B(
        \scalestate_0/PLUSETIME90_m[12] ), .C(
        \scalestate_0/S_DUMPTIME_m[12] ), .Y(
        \scalestate_0/timecount_20_iv_6[12] ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_14  (.A(
        \top_code_0_sigtimedata[3] ), .B(
        \ClockManagement_0/long_timer_0/count[3]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_3 ));
    MX2 \scalestate_0/strippluse_RNO_2[1]  (.A(
        \scalestate_0/STRIPNUM180_NUM[1]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[1]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_421 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m69  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_70 ));
    DFN1 \scalestate_0/strippluse[10]  (.D(
        \scalestate_0/strippluse_RNO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[10] ));
    NOR2A \state_1ms_0/timecount_RNO_5[2]  (.A(
        \state_1ms_0/CS[5]_net_1 ), .B(
        \state_1ms_0/PLUSETIME[2]_net_1 ), .Y(
        \state_1ms_0/PLUSETIME_i_m[2] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m262  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_261 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_262 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_263 ));
    NOR2A \scalestate_0/timecount_ret_85_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[11]_net_1 ), .B(\scalestate_0/N_1089 )
        , .Y(\scalestate_0/S_DUMPTIME_m[11] ));
    DFN1 \PLUSE_0/qq_coder_0/i[2]  (.D(\PLUSE_0/qq_coder_0/i_RNO_2[2] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_4[2] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m76  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_77 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_15_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net )
        , .C(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_20_net ), 
        .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_14_net ));
    NOR3A \top_code_0/relay_close_1_sqmuxa_0_a2_0_0  (.A(
        \top_code_0/N_337 ), .B(\top_code_0/N_154 ), .C(
        \top_code_0/N_147 ), .Y(
        \top_code_0/relay_close_1_sqmuxa_0_a2_0_net_1 ));
    DFN1 \scalestate_0/necount[0]  (.D(
        \scalestate_0/necount_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[0]_net_1 ));
    DFN1 \timer_top_0/timer_0/timedata[16]  (.D(
        \timer_top_0/timer_0/timedata_4[16] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[16]_net_1 ));
    DFN1 \scalestate_0/necount[2]  (.D(
        \scalestate_0/necount_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[2]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[8]  (.D(
        \DUMP_0/dump_coder_0/para4_4[8]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[8]_net_1 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_2_RNO  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0_0 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[2]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0 )
        );
    AO1A \DDS_0/dds_state_0/para_RNO_2[30]  (.A(
        \top_code_0_dds_configdata[13] ), .B(\DDS_0/dds_state_0/N_569 )
        , .C(\DDS_0/dds_state_0/N_514 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[30] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_52_i ));
    DFN1 \top_code_0/scale_rst_2  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_2));
    DFN1E1 \scalestate_0/timecount_ret  (.D(
        \scalestate_0/timecount_cnst[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_cnst_reto[5] ));
    DFN1E1 \scalestate_0/CUTTIME180[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[13]_net_1 )
        );
    DFN1E1 \ClockManagement_0/long_timer_0/count[5]  (.D(
        \ClockManagement_0/long_timer_0/count_n5 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[5]_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[2]  (.D(
        \top_code_0_dds_configdata[1] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[2]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[7] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_3_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ));
    XO1 \PLUSE_0/qq_coder_1/i_reg10_NE_0[0]  (.A(\PLUSE_0/count_7[4] ), 
        .B(\PLUSE_0/qq_para3[4] ), .C(\PLUSE_0/qq_para3[5] ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_NE_0[0]_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[12]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[12] ));
    DFN1 \DUMP_OFF_1/off_on_state_0/cs[1]  (.D(
        \DUMP_OFF_1/off_on_state_0/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/off_on_state_0/cs[1]_net_1 ));
    OA1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO[12]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_208 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[12]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[12]_net_1 ));
    DFN1E1 \scalestate_0/NE_NUM[0]  (.D(\top_code_0_scaledatain[0] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[0]_net_1 ));
    DFN1E1 \plusestate_0/timecount_1[2]  (.D(
        \plusestate_0/timecount_5[2] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[2] ));
    DFN1E1 \top_code_0/pd_pluse_load  (.D(\top_code_0/N_82 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pd_pluse_load));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_21  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_69_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_141_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_21_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_18[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[19]_net_1 ), .B(
        \sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_19[0] ));
    MX2B \plusestate_0/timecount_1_RNO[7]  (.A(\plusestate_0/N_78 ), 
        .B(\plusestate_0/N_253 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[7] ));
    DFN1E0 \DDS_0/dds_state_0/para[30]  (.D(\DDS_0/dds_state_0/N_169 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[30]_net_1 ));
    AO18 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m17  (.A(
        \top_code_0_n_divnum_0[8] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i4_mux ), .C(
        \top_code_0_n_divnum_0[3] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i6_mux ));
    MX2 \plusestate_0/timecount_1_RNO_0[8]  (.A(
        \plusestate_0/DUMPTIME[8]_net_1 ), .B(
        \plusestate_0/PLUSETIME[8]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_79 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[9]_net_1 ));
    AO1 \scalestate_0/timecount_ret_56_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[19]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[19] ), .Y(
        \scalestate_0/timecount_20_0_iv_2[19] ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_0  (.A(
        \scalestate_0/NE_NUM[3]_net_1 ), .B(
        \scalestate_0/necount[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_0_Y ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[4]  (.A(
        \ClockManagement_0/long_timer_0/count_c3 ), .B(
        \ClockManagement_0/long_timer_0/count[4]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n4 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[16]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[16]_net_1 )
        );
    OR2B \plusestate_0/timecount_1_RNO_1[8]  (.A(
        \plusestate_0/CS[8]_net_1 ), .B(top_code_0_pluse_rst), .Y(
        \plusestate_0/N_215 ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[8]  (.A(\scalestate_0/N_555 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[8]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_95  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_95_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_99  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_99_Y ));
    DFN1E1 \scalestate_0/PLUSETIME180[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[10]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m283  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_284 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[0]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/un1_noise_addr_0_i[0] )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ));
    NOR2B \scalestate_0/timecount_ret_11_RNO_3  (.A(
        \scalestate_0/OPENTIME[7]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[7] ));
    XO1 \DUMP_0/dump_coder_0/para6_RNISIH91[2]  (.A(
        \DUMP_0/count_1[2] ), .B(\DUMP_0/dump_coder_0/para6[2]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/i_reg16_1[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_3[0] ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[9]  (.A(
        \top_code_0_dumpdata_0[9] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[9] ));
    DFN1 \ClockManagement_0/long_timer_0/timeup  (.D(
        \ClockManagement_0/long_timer_0/timeup_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(sigtimeup_c));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3_I_9  (
        .A(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/N_2 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNILKJB2[3]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[3] ));
    DFN1 \top_code_0/scale_start_ret_2  (.D(\xa_c[0] ), .CLK(GLA_net_1)
        , .Q(\top_code_0/xa_c_reto[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_152  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_102_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_65_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_152_Y ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_17  (.A(
        \timer_top_0/dataout[17] ), .B(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_17_Y ));
    NOR2B \DUMP_0/dump_state_0/cs_RNIBSCA[3]  (.A(
        \DUMP_0/dump_state_0/cs[3]_net_1 ), .B(\DUMP_0/i_2[1] ), .Y(
        \DUMP_0/dump_state_0/N_195 ));
    NOR2 \top_code_0/state_1ms_lc_1_sqmuxa_0_a2_0  (.A(
        \top_code_0/N_157 ), .B(\top_code_0/N_163 ), .Y(
        \top_code_0/state_1ms_lc_1_sqmuxa_0_a2_0_net_1 ));
    NOR2A \scalestate_0/strippluse_RNO_1[3]  (.A(\scalestate_0/N_423 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[3] ));
    NOR2B \sd_acq_top_0/sd_sacq_state_0/cs4_0_o2  (.A(
        \sd_acq_top_0/i_10[0] ), .B(net_27), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ));
    NOR2A \scalestate_0/timecount_ret_0_RNIT4EE  (.A(
        \scalestate_0/timecount_cnst_m_0_reto[6] ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .Y(
        \scalestate_0/timecount_cnst_m_reto[6] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m29  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_28 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_29 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_30 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_16  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[1] )
        , .C(\s_acq_change_0_s_stripnum[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8 ));
    NOR3B \plusestate_0/soft_d_RNO_1  (.A(\plusestate_0/N_302 ), .B(
        \plusestate_0/N_301 ), .C(\plusestate_0/CS[5]_net_1 ), .Y(
        \plusestate_0/N_299 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m240  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_239 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_240 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_241 ));
    DFN1E1 \top_code_0/noisedata[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[9] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[8] ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m44_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[3]_net_1 ));
    DFN1 \DUMP_OFF_0/off_on_timer_0/count[2]  (.D(
        \DUMP_OFF_0/off_on_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/count_3[2] ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_4  (.A(
        \scalestate_0/necount_cmp_0/NOR3A_2_Y ), .B(
        \scalestate_0/necount_cmp_0/OR2A_4_Y ), .C(
        \scalestate_0/necount_cmp_0/NAND3A_5_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_4_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_7_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_9_net ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[9] ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_net_1 ));
    AO1 \DDS_0/dds_state_0/para_RNO_2[7]  (.A(
        \DDS_0/dds_state_0/para[7]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569 ), .C(\DDS_0/dds_state_0/N_270 ), .Y(
        \DDS_0/dds_state_0/para_9_i_i_1[7] ));
    DFN1E1 \top_code_0/s_addchoice[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice[4] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_9  (.A(\xd_in[5] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[5] ));
    DFN1 \scalestate_0/CS[14]  (.D(\scalestate_0/CS_RNO[14]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[14]_net_1 ));
    AO1 \noisestate_0/dumpoff_ctr_RNO_0  (.A(noisestate_0_dumpoff_ctr), 
        .B(\noisestate_0/N_250 ), .C(\noisestate_0/CS[5]_net_1 ), .Y(
        \noisestate_0/N_112 ));
    NOR2A \state_1ms_0/timecount_RNO_6[5]  (.A(
        \state_1ms_0/CS[8]_net_1 ), .B(\state_1ms_0/CUTTIME[5]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_i_m[5] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i4_mux ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[6]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[6] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[6]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m143  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_128 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_143 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[3] ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[15]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_245 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO[15]_net_1 ));
    DFN1C0 \bridge_div_0/count[2]  (.D(\bridge_div_0/count_5[2] ), 
        .CLK(ddsclkout_c), .CLR(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[2]_net_1 ));
    MX2 \top_code_0/state_1ms_start_ret_2_RNIPLG71  (.A(
        \top_code_0/top_code_0_state_1ms_start_reto ), .B(
        \top_code_0/un1_xa_4_reto ), .S(\top_code_0/N_112_reto ), .Y(
        \top_code_0/N_795_reto ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[6]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[6] ));
    DFN1E1 \noisestate_0/timecount_1[9]  (.D(
        \noisestate_0/timecount_5[9] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[9] ));
    DFN1E1 \top_code_0/plusedata[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[2] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[14]  (.A(
        \DDS_0/dds_state_0/para[14]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_461 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[14] ));
    NOR3C \DUMP_OFF_1/off_on_coder_0/i_RNO[1]  (.A(
        nsctrl_choice_0_dumponoff_rst), .B(
        \DUMP_OFF_1/off_on_coder_0/i_0_1[1] ), .C(
        \DUMP_OFF_1/off_on_coder_0/i_0_2[1] ), .Y(
        \DUMP_OFF_1/off_on_coder_0/i_RNO_4[1] ));
    DFN1E1 \top_code_0/bri_datain[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[5] ));
    DFN1E1 \scalestate_0/PLUSETIME90[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[15]_net_1 ));
    DFN1 \top_code_0/relay_close[9]  (.D(
        \top_code_0/relay_close_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[9] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m126  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_123 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_126 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_127 ));
    NOR2B \ClockManagement_0/clk_10k_0/un1_count_1_I_44  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_TMP[0] ), .B(
        \ClockManagement_0/clk_10k_0/count[1]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_1[0] ));
    NOR2A \scanstate_0/timecount_1_RNO[1]  (.A(\scanstate_0/N_59 ), .B(
        \scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[1] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[11]_net_1 ));
    DFN1E1 \top_code_0/change[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/change_1_sqmuxa ), .Q(
        \top_code_0_change[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[11]  (.D(
        \DUMP_0/dump_coder_0/para5_4[11] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[11]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i16_mux ));
    DFN1 \DUMP_0/dump_state_0/cs_i_0[0]  (.D(\DUMP_0/dump_state_0/cs4 )
        , .CLK(GLA_net_1), .Q(\DUMP_0/dump_state_0/cs_i_0[0]_net_1 ));
    NOR2 \scalestate_0/CS_RNIKSD4[19]  (.A(\scalestate_0/CS[19]_net_1 )
        , .B(\scalestate_0/CS[20]_net_1 ), .Y(\scalestate_0/N_1262 ));
    DFN1E1 \noisestate_0/acqtime[15]  (.D(\top_code_0_noisedata[15] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[15]_net_1 ));
    DFN1 \CAL_0/cal_div_0/count[1]  (.D(\CAL_0/cal_div_0/count_5[1] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[1]_net_1 ));
    MX2 \top_code_0/relay_on_RNO_0[3]  (.A(\relay_on_c[3] ), .B(
        \GPMI_0_dataout[3] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_812 ));
    DFN1E1 \scalestate_0/timecount[21]  (.D(
        \scalestate_0/timecount_20[21] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(\scalestate_0_timecount[21] ));
    OA1B \state_1ms_0/CS_RNO[4]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[4] ), 
        .Y(\state_1ms_0/CS_RNO_3[4] ));
    OR3 \state_1ms_0/timecount_RNO_1[13]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[13] ), .B(
        \state_1ms_0/CUTTIME_m[13] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[13] ), .Y(
        \state_1ms_0/timecount_8[13] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m295  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_296 ));
    NOR2B \bri_dump_sw_0/dumpoff_ctr_RNO  (.A(
        \bri_dump_sw_0/dumpoff_ctr_5 ), .B(net_27), .Y(
        \bri_dump_sw_0/dumpoff_ctr_RNO_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[13]_net_1 ));
    MX2 \n_acq_change_0/n_rst_n_5  (.A(top_code_0_pluse_rst_0), .B(
        top_code_0_noise_rst_0), .S(top_code_0_pluse_noise_ctrl), .Y(
        \n_acq_change_0/n_rst_n_5_net_1 ));
    OA1B \top_code_0/pluseload_RNO  (.A(\top_code_0/N_164 ), .B(
        \top_code_0/N_175 ), .C(\top_code_0/N_297 ), .Y(
        \top_code_0/N_90 ));
    DFN1 \GPMI_0/xwe_xzcs2_syn_0/code_en  (.D(
        \GPMI_0/xwe_xzcs2_syn_0/code_en_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(GPMI_0_code_en));
    NOR2B \ClockManagement_0/long_timer_0/count_RNI8RES3[8]  (.A(
        \ClockManagement_0/long_timer_0/count_c7 ), .B(
        \ClockManagement_0/long_timer_0/count[8]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c8 ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_1_i_a2_0  
        (.A(\top_code_0_sd_sacq_choice[3] ), .B(
        \top_code_0_sd_sacq_choice[1] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_1_i_a2_0_net_1 )
        );
    NOR3C \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa  (.A(OR2_1_Y), .B(
        \DUMP_ON_0/off_on_state_0_state_over ), .C(OR2_2_Y), .Y(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ));
    DFN1 \scalestate_0/CS[11]  (.D(\scalestate_0/CS_RNIRUEO[10]_net_1 )
        , .CLK(GLA_net_1), .Q(\scalestate_0/CS[11]_net_1 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_5_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(\pd_pluse_top_0/count_6[3] ), .C(
        \pd_pluse_top_0/count_6[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_5_net ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_46  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_78_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_31_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_46_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[7]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI4G0P[14]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[14]_net_1 ), .B(
        \sd_acq_top_0/count_0[14] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_14[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[8]  (.A(
        \state_1ms_0_timecount[8] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_247 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[10]  (.D(
        \DUMP_0/dump_coder_0/para4_4[10]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[10]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[20]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[20]_net_1 ));
    DFN1 \DUMP_0/off_on_coder_0/i[1]  (.D(
        \DUMP_0/off_on_coder_0/i_RNO_2[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_0[1] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_56_i ));
    XO1 \scalestate_0/fst_lst_pulse_RNO_8  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/NE_NUM[6]_net_1 ), .C(
        \scalestate_0/fst_lst_pulse8_5 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_1 ));
    NOR3C \DUMP_0/off_on_coder_0/i_RNO[1]  (.A(
        \DUMP_0/off_on_coder_0/i_0_2[1] ), .B(
        \DUMP_0/off_on_coder_0/i_0_1[1] ), .C(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_coder_0/i_RNO_2[1] ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_4  (.A(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .B(
        \timer_top_0/dataout[21] ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_10_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_4_Y ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[8] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_56_i ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m44_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[15] ));
    DFN1E1 \plusestate_0/DUMPTIME[13]  (.D(\top_code_0_plusedata[13] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[13]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m70  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m70_0 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_34  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_161_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_108_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_34_Y ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_8  
        (.A(\s_acq_change_0_s_stripnum[0] ), .B(
        \s_acq_change_0_s_stripnum[1] ), .C(
        \s_acq_change_0_s_stripnum[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11 ));
    DFN1 \timer_top_0/state_switch_0/clk_en_pluse  (.D(
        \timer_top_0/state_switch_0/clk_en_pluse_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(timer_top_0_clk_en_pluse));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_54_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[0] )
        );
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIG6DM[7]  (.A(
        \sd_acq_top_0/count_3[7] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[7]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_5[0] ));
    DFN1 \DDS_0/dds_timer_0/count[6]  (.D(\DDS_0/dds_timer_0/count_n6 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[6] ));
    OA1 \scalestate_0/CS_i_RNO[0]  (.A(timer_top_0_clk_en_scale_0), .B(
        \scalestate_0/CS_i[0]_net_1 ), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/CS_i_RNO_0[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[0]  (.D(
        \DUMP_0/dump_coder_0/para2_4[0]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[0]_net_1 ));
    DFN1E1 \top_code_0/sigtimedata[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[10] ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/data[1]  (.D(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[1]_net_1 ), .CLK(
        GLA_net_1), .Q(\DSTimer_0/dump_sustain_timer_0/data[1]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_47_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[16]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[16] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_16[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[11]_net_1 ), 
        .B(\pd_pluse_top_0/count_0[11] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_11[0] ));
    AOI1 \scalestate_0/necount_cmp_0/AOI1_ALEB  (.A(
        \scalestate_0/necount_cmp_0/AND3_0_Y ), .B(
        \scalestate_0/necount_cmp_0/AO1_1_Y ), .C(
        \scalestate_0/necount_cmp_0/AO1_0_Y ), .Y(
        \scalestate_0/necount_LE_M_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_54_i ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[21]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[21]_net_1 ));
    XOR2 \PLUSE_0/qq_coder_1/un1_qq_para2_0[0]  (.A(
        \PLUSE_0/qq_para2[0] ), .B(\PLUSE_0/count_7[0] ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_0[0]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[7]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[7] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_RNO  (
        .A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop ), 
        .B(scan_scale_sw_0_s_start), .C(
        \Signal_Noise_Acq_0/signal_acq_0/clkout ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_4 ));
    AO1 \scalestate_0/timecount_ret_25_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL[11]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[11] )
        , .Y(\scalestate_0/timecount_20_iv_3[11] ));
    MX2 \scalestate_0/CS_RNO_0[15]  (.A(\scalestate_0/CS[15]_net_1 ), 
        .B(\scalestate_0/CS[14]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1228 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[14]  (.A(
        \s_acq_change_0/s_acqnum_5[14] ), .B(
        \s_acq_change_0_s_acqnum[14] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_84 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[2]  (.A(
        \scanstate_0_timecount[2] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_231 ));
    DFN1E1 \scanstate_0/dectime[12]  (.D(\top_code_0_scandata[12] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[12]_net_1 ));
    DFN1 \DDS_0/dds_state_0/fq_ud_reg  (.D(
        \DDS_0/dds_state_0/fq_ud_reg_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/fq_ud_reg_net_1 ));
    DFN1E1 \top_code_0/pd_pluse_choice[3]  (.D(\GPMI_0_dataout[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_choice_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_choice[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m42_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[17] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[3]  (.D(
        \DUMP_0/dump_coder_0/para5_4[3] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[3]_net_1 ));
    DFN1E1 \top_code_0/bri_datain[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[4] ));
    XOR3 \bridge_div_0/dataall_1_I_14  (.A(\top_code_0_scaleddsdiv[2] )
        , .B(\top_code_0_scaleddsdiv[5] ), .C(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_1[0] ), .Y(
        \bridge_div_0/dataall_1[2] ));
    IOTRI_OB_EB \calcuinter_pad/U0/U1  (.D(calcuinter_c), .E(VCC), 
        .DOUT(\calcuinter_pad/U0/NET1 ), .EOUT(
        \calcuinter_pad/U0/NET2 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[7]  (.D(\top_code_0_scaledatain[7] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[7]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[10] ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/HOR2_10_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_13_net ), 
        .B(\pd_pluse_top_0/count[13] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[13] ));
    XOR3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m13  (.A(
        \top_code_0_n_divnum_0[1] ), .B(\top_code_0_n_divnum_0[6] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_i ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_14_i ));
    DFN1E1 \top_code_0/n_divnum[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[4] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m47_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[10]  (.D(
        \top_code_0_pd_pluse_data[10] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[10]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[17]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[17]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_499 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/signal_data_t_0_11  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] ), .Y(
        \Signal_Noise_Acq_0/un1_signal_acq_0[3] ));
    DFN1 \DUMP_ON_0/off_on_timer_0/count[0]  (.D(
        \DUMP_ON_0/off_on_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/count_5[0] ));
    IOPAD_TRI \ddsreset_pad/U0/U0  (.D(\ddsreset_pad/U0/NET1 ), .E(
        \ddsreset_pad/U0/NET2 ), .PAD(ddsreset));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_34  (.A(
        \ClockManagement_0/clk_10k_0/count[6]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_11[0] ), 
        .Y(\ClockManagement_0/clk_10k_0/I_34_0 ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_70_i ));
    IOPAD_IN \xa_pad[7]/U0/U0  (.PAD(xa[7]), .Y(\xa_pad[7]/U0/NET1 ));
    OR2A \topctrlchange_0/sw_acq1_RNO  (.A(net_27), .B(
        \topctrlchange_0/N_10 ), .Y(
        \topctrlchange_0/sw_acq1_RNO_1_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME90[8]  (.D(\top_code_0_scaledatain[8] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[8]_net_1 ));
    OAI1 \scalestate_0/CS_RNI59HI[4]  (.A(\scalestate_0/CS[10]_net_1 ), 
        .B(\scalestate_0/CS[4]_net_1 ), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/N_1093 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m19  
        (.A(\s_acq_change_0_s_stripnum[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[6]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i12_mux )
        );
    XOR2 \DUMP_0/dump_coder_0/para3_RNIEJFH[3]  (.A(
        \DUMP_0/dump_coder_0/para3[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_3[0] ));
    NOR2B \state_1ms_0/timecount_RNO_1[18]  (.A(
        \state_1ms_0/CUTTIME[18]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/timecount_8[18] ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_6  (.A(\ADC_c[4] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_6 ));
    NOR2B \scalestate_0/timecount_ret_41_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[2]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[2] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_14_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_14_net ));
    IOPAD_IN \ADC_pad[9]/U0/U0  (.PAD(ADC[9]), .Y(\ADC_pad[9]/U0/NET1 )
        );
    DFN1 \noisestate_0/rt_sw  (.D(\noisestate_0/rt_sw_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(noisestate_0_rt_sw));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[1] ), .CLK(
        GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_25_RNO_0  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[11]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[11] ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_8  (.A(\ADC_c[2] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_8 ));
    NOR2A \top_code_0/noise_start_ret_3_RNO_0  (.A(\top_code_0/N_332 ), 
        .B(\top_code_0/N_149 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_44_i_a2_0 ));
    AND2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_31  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[5] ));
    DFN1 \DUMP_0/dump_state_0/cs[6]  (.D(
        \DUMP_0/dump_state_0/cs_nsss[6] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[6]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_7  (.A(\ADC_c[3] ), 
        .B(top_code_0_n_s_ctrl), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]  (
        .D(\top_code_0_n_acqnum_2[10] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]_net_1 )
        );
    IOBI_IB_OB_EB \xd_pad[5]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[5] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[5]/U0/NET3 ), .DOUT(\xd_pad[5]/U0/NET1 ), .EOUT(
        \xd_pad[5]/U0/NET2 ), .Y(\xd_in[5] ));
    NOR3A \top_code_0/un1_xa_8_16_i_i_o3_i_a2_5  (.A(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_3_net_1 ), .B(\xa_c[14] ), 
        .C(\xa_c[15] ), .Y(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_5_net_1 ));
    DFN1E1 \top_code_0/cal_load  (.D(\top_code_0/N_64 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_cal_load));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m46  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_47 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[6]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNIOEM12[4]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c2 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c4 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[4]  (.D(
        \DUMP_0/dump_coder_0/para4_4[4]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[4]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_3[4]  (.A(
        \state_1ms_0/CUTTIME[4]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[4] ));
    XA1 \PLUSE_0/qq_timer_0/count_RNO[2]  (.A(
        \PLUSE_0/qq_timer_0/count_c1 ), .B(\PLUSE_0/count_9[2] ), .C(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_0/count_n2 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_0  (.A(
        \timer_top_0/dataout[16] ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_7_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_0_Y ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[7]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[7] ));
    AND2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_8_inst  (.A(
        \sd_acq_top_0/count_3[6] ), .B(\sd_acq_top_0/count_3[7] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_8_net ));
    NOR2B \scalestate_0/CS_RNO[10]  (.A(\scalestate_0/N_1224 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO[10]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[3]  (.D(
        \DUMP_0/dump_coder_0/para2_4[3]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_48  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_113_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_136_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_48_Y ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_11  (.A(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .B(
        \timer_top_0/dataout[17] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_11_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[2] ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/start  (.D(
        \DSTimer_0/dump_sustain_timer_0/start11 ), .CLK(clock_10khz), 
        .Q(net_40));
    AX1C \ClockManagement_0/clk_10k_0/un1_count_1_I_36  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_11[0] ), 
        .B(\ClockManagement_0/clk_10k_0/count[6]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/I_36_0 ));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[6]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_186 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_185 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[6]_net_1 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_32  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m39 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[8] )
        );
    NOR2B \state_1ms_0/timecount_RNO[19]  (.A(\state_1ms_0/N_86 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[19]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[4]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[4] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_2[4] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[10]  (.D(
        \top_code_0_pd_pluse_data[10] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[10]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[11]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[11] ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/signal_data_t_0_14  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] ), .Y(
        \Signal_Noise_Acq_0/un1_signal_acq_0[0] ));
    XOR2 \bridge_div_0/count_5_I_9  (.A(\bridge_div_0/N_4 ), .B(
        \bridge_div_0/count_RNIHPOM7[3]_net_1 ), .Y(
        \bridge_div_0/count_5[3] ));
    NOR2A \scalestate_0/timecount_ret_67_RNO_0  (.A(
        \scalestate_0/ACQTIME[14]_net_1 ), .B(\scalestate_0/N_1065 ), 
        .Y(\scalestate_0/ACQTIME_m[14] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[5]  (.A(
        \scalestate_0/s_acqnum_7[5] ), .B(\scalestate_0_s_acqnum[5] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_552 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_1_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        );
    IOBI_IB_OB_EB \xd_pad[0]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[0] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[0]/U0/NET3 ), .DOUT(\xd_pad[0]/U0/NET1 ), .EOUT(
        \xd_pad[0]/U0/NET2 ), .Y(\xd_in[0] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[3]  (.D(
        \top_code_0_n_acqnum_2[3] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[3]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[4] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[0] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNITTM5[3]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[3]_net_1 ), .B(
        \sd_acq_top_0/count_10[3] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_3[0] ));
    DFN1 \scanstate_0/dumpoff_ctr  (.D(\scanstate_0/dumpoff_ctr_RNO_3 )
        , .CLK(GLA_net_1), .Q(scanstate_0_dumpoff_ctr));
    NOR3C \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa  (.A(
        \DUMP_OFF_0/off_on_state_0_state_over ), .B(
        bri_dump_sw_0_dumpoff_ctr), .C(bri_dump_sw_0_reset_out), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ));
    OR3A \scalestate_0/intertodsp_RNO_1  (.A(\scalestate_0/N_1196 ), 
        .B(\scalestate_0/un1_CS_27 ), .C(
        \scalestate_0/intertodsp_1_sqmuxa ), .Y(
        \scalestate_0/un1_CS6_14 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m279  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_272 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_279 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[14] ));
    DFN1 \DUMP_0/off_on_coder_1/i[1]  (.D(
        \DUMP_0/off_on_coder_1/i_RNO_1[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_1[1] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[5] ));
    DFN1E1 \scalestate_0/OPENTIME[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[11]_net_1 ));
    IOPAD_TRI \relay_close_pad[7]/U0/U0  (.D(
        \relay_close_pad[7]/U0/NET1 ), .E(\relay_close_pad[7]/U0/NET2 )
        , .PAD(relay_close[7]));
    DFN1 \DDS_0/dds_coder_0/i[1]  (.D(
        \DDS_0/dds_coder_0/i_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/i[1] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[2]  (.A(
        \top_code_0_s_acqnum_2[2] ), .B(\scalestate_0_s_acqnum[2] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[2] ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[6]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[6]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/i_0[6] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[10]_net_1 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[10]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[10]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m232  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_231 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_232 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_233 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ));
    AO1 \scalestate_0/timecount_ret_28_RNO_6  (.A(
        \scalestate_0/CUTTIME180_TEL[1]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[1] ), 
        .Y(\scalestate_0/timecount_20_iv_3[1] ));
    NOR3C \DUMP_0/dump_coder_0/i_RNO_1[3]  (.A(
        \DUMP_0/dump_coder_0/i_0_0_a2_7[3] ), .B(
        \DUMP_0/dump_coder_0/i_0_0_a2_6[3] ), .C(
        \DUMP_0/dump_coder_0/i_0_0_a2_8[3] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_10[3] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m73  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_72 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_73 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_74 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[4] ));
    AO1A \scalestate_0/timecount_ret_13_RNIQQ31  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .B(
        \scalestate_0/timecount_cnst_m_0_reto[9] ), .C(
        \scalestate_0/timecount_20_iv_10_reto[9] ), .Y(
        \scalestate_0_timecount[9] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[9]  (.A(
        \scalestate_0/s_acqnum_7[9] ), .B(\scalestate_0_s_acqnum[9] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_556 ));
    DFN1 \DUMP_0/off_on_coder_0/i[0]  (.D(
        \DUMP_0/off_on_coder_0/i_RNO_2[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_0[0] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i18_mux ));
    NOR2B \scalestate_0/strippluse_RNO[9]  (.A(\scalestate_0/N_568 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[9]_net_1 ));
    AO1A \topctrlchange_0/sw_acq1_RNO_1  (.A(scalestate_0_sw_acq1), .B(
        \top_code_0_change_0[0] ), .C(\topctrlchange_0/sw_acq1in3_i_m )
        , .Y(\topctrlchange_0/sw_acq1_6_iv ));
    NOR3C \scalestate_0/timecount_ret_61_RNO_1  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[12]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[12] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[4]  (.D(
        \top_code_0_halfdata_0[4] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[4] ));
    OA1 \noisestate_0/CS_i_0_RNO[0]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS_li[0] ), .C(top_code_0_noise_rst), .Y(
        \noisestate_0/CS_i_0_RNO[0]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m41_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[18] ));
    NOR3B \scalestate_0/M_pulse_RNIJJN9  (.A(
        \scalestate_0/M_pulse_net_1 ), .B(\scalestate_0/CS[15]_net_1 ), 
        .C(\scalestate_0/necount_LE_M_net_1 ), .Y(
        \scalestate_0/timecount_16_sqmuxa_1 ));
    IOTRI_OB_EB \relay_on_pad[8]/U0/U1  (.D(\relay_on_c[8] ), .E(VCC), 
        .DOUT(\relay_on_pad[8]/U0/NET1 ), .EOUT(
        \relay_on_pad[8]/U0/NET2 ));
    NOR2 \DUMP_OFF_0/off_on_coder_0/i_RNO_1[1]  (.A(
        \DUMP_OFF_0/count_3[1] ), .B(\DUMP_OFF_0/count_3[0] ), .Y(
        \DUMP_OFF_0/off_on_coder_0/i_0_1[1] ));
    DFN1 \DUMP_0/off_on_timer_0/count[2]  (.D(
        \DUMP_0/off_on_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_2[2] ));
    DFN1E1 \top_code_0/s_periodnum[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_periodnum_1_sqmuxa ), .Q(
        \top_code_0_s_periodnum[1] ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[10]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[10]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/i[10] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIE04O4[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_3[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_2[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_17[0] ));
    NOR2A \scalestate_0/timecount_ret_35_RNO_4  (.A(
        \scalestate_0/ACQTIME[9]_net_1 ), .B(\scalestate_0/N_1065 ), 
        .Y(\scalestate_0/ACQTIME_m[9] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_8  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_8_Y ));
    AO1C \plusestate_0/dds_config_RNO_0  (.A(
        \plusestate_0/CS[9]_net_1 ), .B(plusestate_0_dds_config), .C(
        \plusestate_0/N_301 ), .Y(\plusestate_0/N_142 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para1[0]  (.D(
        \top_code_0_bri_datain[0] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para1[0] ));
    NOR2B \state_1ms_0/reset_out_RNO  (.A(\state_1ms_0/N_154 ), .B(
        top_code_0_state_1ms_rst_n), .Y(\state_1ms_0/reset_out_RNO_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m43_6 ));
    NOR2B \PLUSE_0/qq_timer_0/count_RNO_0[4]  (.A(\PLUSE_0/count_9[3] )
        , .B(\PLUSE_0/qq_timer_0/count_c2 ), .Y(
        \PLUSE_0/qq_timer_0/count_9_0 ));
    NOR2B \state_1ms_0/timecount_RNO[6]  (.A(\state_1ms_0/N_73 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[6]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNIH9JE  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_net_1 ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/clk_add_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_80  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_80_Y ));
    AO1C \noisestate_0/CS_RNO_0[3]  (.A(\noisestate_0/CS[2]_net_1 ), 
        .B(timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[3] ));
    DFN1 \PLUSE_0/qq_coder_0/i[1]  (.D(\PLUSE_0/qq_coder_0/i_RNO_6[1] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_9[1] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[2]  (.D(
        \top_code_0_halfdata_0[2] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[2] ));
    OR3 \scalestate_0/timecount_ret_47_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[16] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[16] ), .C(
        \scalestate_0/timecount_20_0_iv_2[16] ), .Y(
        \scalestate_0/timecount_20_0_iv_4[16] ));
    NOR3B \scalestate_0/CUTTIMEI90_538_e  (.A(\scalestate_0/N_64 ), .B(
        \scalestate_0/N_65 ), .C(\top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/N_1751 ));
    IOPAD_IN \xa_pad[1]/U0/U0  (.PAD(xa[1]), .Y(\xa_pad[1]/U0/NET1 ));
    NOR3C \GPMI_0/xwe_xzcs2_syn_0/code_en_RNO  (.A(
        \GPMI_0/xwe_xzcs2_syn_0/code_en_0_0 ), .B(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_net_1 ), .C(net_27), .Y(
        \GPMI_0/xwe_xzcs2_syn_0/code_en_RNO_net_1 ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_10_RNO  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_10_0 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_8 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_5 )
        );
    NOR2A \scanstate_0/timecount_1_RNO[15]  (.A(\scanstate_0/N_73 ), 
        .B(\scanstate_0/N_233 ), .Y(\scanstate_0/timecount_5[15] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[5]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[5] ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIG6I21[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_12_0 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_3 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_2 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m12  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_13_0 ));
    DFN1E1 \scalestate_0/ACQTIME[12]  (.D(\top_code_0_scaledatain[12] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[12]_net_1 ));
    AX1C \DDS_0/dds_timer_0/count_RNO_0[6]  (.A(\DDS_0/count[5] ), .B(
        \DDS_0/dds_timer_0/count_c4 ), .C(\DDS_0/count[6] ), .Y(
        \DDS_0/dds_timer_0/count_n6_tz ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI68EB[5]  (.A(
        \sd_acq_top_0/count_3[5] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[5]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_7[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_1[0] ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2b_9_inst  
        (.A(\pd_pluse_top_0/count_6[0] ), .B(
        \pd_pluse_top_0/count_6[1] ), .C(\pd_pluse_top_0/count_6[2] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net )
        );
    NOR2B \noisestate_0/acqtime_0_sqmuxa  (.A(top_code_0_nstatechoice), 
        .B(top_code_0_nstateload), .Y(
        \noisestate_0/acqtime_0_sqmuxa_net_1 ));
    DFN1P0 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]  
        (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[0]_net_1 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .PRE(
        s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        );
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[5]_net_1 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[12]_net_1 ));
    XA1C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_17[4]  (.A(
        \pd_pluse_top_0/count_1[5] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[5]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_2[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_4[4] ));
    OA1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_20  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_6 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_7 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_11 ));
    DFN1 \CAL_0/cal_div_0/count[4]  (.D(\CAL_0/cal_div_0/count_5[4] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[4]_net_1 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_10_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net ), 
        .B(\pd_pluse_top_0/count_0[9] ), .C(
        \pd_pluse_top_0/count_0[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_14_net ));
    DFN1E1 \state_1ms_0/CUTTIME[14]  (.D(
        \top_code_0_state_1ms_data[14] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[14]_net_1 ));
    AO1 \PLUSE_0/bri_coder_0/half_0_I_25  (.A(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[1] ), .B(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[2] ), .C(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[0] ), .Y(
        \PLUSE_0/bri_coder_0_half ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_3_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_3_net ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[7]  (.A(
        \top_code_0_dumpdata_0[7] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[7] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_55  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_55_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_59  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_59_Y ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNI7UUI2[5]  (.A(
        \ClockManagement_0/long_timer_0/count_c4 ), .B(
        \ClockManagement_0/long_timer_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c5 ));
    DFN1E1 \scalestate_0/timecount_ret_79  (.D(
        \scalestate_0/un1_timecount_2_sqmuxa_9 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/un1_timecount_2_sqmuxa_9_reto ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[5]  (.D(
        \top_code_0_pd_pluse_data[5] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[5]_net_1 ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        );
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[6]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[6] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_1[6] ));
    DFN1E1 \scanstate_0/timecount_1[12]  (.D(
        \scanstate_0/timecount_5[12] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[12] ));
    IOPAD_TRI \relay_on_pad[6]/U0/U0  (.D(\relay_on_pad[6]/U0/NET1 ), 
        .E(\relay_on_pad[6]/U0/NET2 ), .PAD(relay_on[6]));
    DFN1E1 \state_1ms_0/PLUSECYCLE[3]  (.D(
        \top_code_0_state_1ms_data[3] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m125  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_124 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_125 ), .S(
        \top_code_0_s_addchoice_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_126 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[8]_net_1 ));
    AO1C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_15  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_4 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_6 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[9] ));
    MX2 \scalestate_0/dump_sustain_ctrl_RNO_0  (.A(
        \scalestate_0/CS_0[11]_net_1 ), .B(
        scalestate_0_dump_sustain_ctrl), .S(\scalestate_0/N_1183 ), .Y(
        \scalestate_0/N_744 ));
    OR3 \DUMP_0/dump_coder_0/para4_RNI8QQC2[10]  (.A(
        \DUMP_0/dump_coder_0/un1_count_1_10[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_0_0[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_1_NE_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_8[0] ));
    NOR2B \top_code_0/state_1ms_start_ret_1_RNI28QI1  (.A(
        \top_code_0/N_799_reto ), .B(\top_code_0/net_27_reto ), .Y(
        top_code_0_noise_start));
    AO1C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_19  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[10]_net_1 )
        , .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_5 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_10 ));
    OR3 \scalestate_0/timecount_ret_32_RNISA41  (.A(
        \scalestate_0/timecount_20_iv_9_reto[4] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[4] ), .C(
        \scalestate_0/timecount_cnst_m_reto[1] ), .Y(
        \scalestate_0_timecount[4] ));
    NOR2A \scalestate_0/strippluse_RNO_1[2]  (.A(\scalestate_0/N_422 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[2] ));
    NOR2B \state_1ms_0/timecount_RNO[15]  (.A(\state_1ms_0/N_82 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[15]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[22]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[23]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_269 ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_5  (.A(
        \scalestate_0/M_NUM[1]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .C(
        \scalestate_0/necount_cmp_0/OR2A_1_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_5_Y ));
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_3  (.A(
        \scalestate_0/NE_NUM[7]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .C(
        \scalestate_0/necount_cmp_1/OR2A_2_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_3_Y ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[2]  (.A(
        \PLUSE_0/bri_state_0/cs[2]_net_1 ), .B(
        \PLUSE_0/bri_state_0/csse_1_0_a4_0_0 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[2] ));
    NOR2A \topctrlchange_0/sw_acq1_RNO_2  (.A(\top_code_0_change[1] ), 
        .B(plusestate_0_sw_acq1), .Y(\topctrlchange_0/sw_acq1in3_i_m ));
    OR3 \top_code_0/sigrst_RNO_0  (.A(\top_code_0/N_151 ), .B(
        \top_code_0/N_158 ), .C(\top_code_0/N_147 ), .Y(
        \top_code_0/N_209 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[0]_net_1 ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[1]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_33 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[1] ));
    NOR3B \top_code_0/un1_state_1ms_rst_n117_47_i_a3  (.A(\xa_c[7] ), 
        .B(\top_code_0/N_339 ), .C(\top_code_0/N_139 ), .Y(
        \top_code_0/N_330 ));
    NOR3C \timer_top_0/state_switch_0/clk_en_st1ms_RNO  (.A(net_27), 
        .B(\timer_top_0/timer_0_time_up ), .C(
        top_code_0_state_1ms_start), .Y(
        \timer_top_0/state_switch_0/clk_en_st1ms_RNO_net_1 ));
    OR3 \PLUSE_0/bri_state_0/cs_RNI2QTF2[1]  (.A(
        \PLUSE_0/bri_state_0/cs[8]_net_1 ), .B(
        \PLUSE_0/bri_state_0/N_181 ), .C(\PLUSE_0/bri_state_0/N_180 ), 
        .Y(\PLUSE_0/bri_state_0/N_145 ));
    XO1 \DUMP_0/dump_coder_0/para3_RNI6HV21[6]  (.A(
        \DUMP_0/count_0[6] ), .B(\DUMP_0/dump_coder_0/para3[6]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_2_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_1[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[5]  (.D(
        \DUMP_0/dump_coder_0/para4_4[5]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[5]_net_1 ));
    DFN1E0 \DDS_0/dds_state_0/para[23]  (.D(\DDS_0/dds_state_0/N_20 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[23]_net_1 ));
    DFN1 \s_acq_change_0/s_stripnum[0]  (.D(
        \s_acq_change_0/s_stripnum_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[0] ));
    MX2B \ClockManagement_0/clk_10k_0/clock_10khz_RNO_0  (.A(
        clock_10khz), .B(clock_10khz), .S(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/clock_10khz_RNO_0_net_1 ));
    DFN1 \scalestate_0/CS[2]  (.D(\scalestate_0/CS_RNO_1[2] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[2]_net_1 ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_70_i ));
    DFN1 \scalestate_0/sw_acq2  (.D(\scalestate_0/sw_acq2_RNO_1 ), 
        .CLK(GLA_net_1), .Q(scalestate_0_sw_acq2));
    AO18 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m7  (.A(
        \top_code_0_n_divnum_0[7] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i2_mux ), .C(
        \top_code_0_n_divnum_0[2] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i4_mux ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[2]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[2] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[2]_net_1 ));
    DFN1 \DDS_0/dds_state_0/cs[1]  (.D(
        \DDS_0/dds_state_0/cs_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[1]_net_1 ));
    NOR3B \scalestate_0/CUTTIME180_432_e  (.A(\scalestate_0/N_60 ), .B(
        \scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/N_1645 ));
    DFN1 \PLUSE_0/qq_state_0/cs[1]  (.D(
        \PLUSE_0/qq_state_0/cs_RNO_1[1] ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_0/cs[1]_net_1 ));
    DFN1E1 \state_1ms_0/PLUSETIME[7]  (.D(
        \top_code_0_state_1ms_data[7] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[7]_net_1 ));
    DFN1E1 \noisestate_0/timecount_1[11]  (.D(
        \noisestate_0/timecount_5[11] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[11] ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_70_i ));
    DFN1E1 \scalestate_0/timecount_ret_55  (.D(
        \scalestate_0/OPENTIME_TEL_m[19] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/OPENTIME_TEL_m_reto[19] ));
    DFN1E1 \noisestate_0/acqtime[12]  (.D(\top_code_0_noisedata[12] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[12]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_9_i_0_a2_4[22]  (.A(\DDS_0/i[0] ), 
        .B(top_code_0_dds_load), .Y(\DDS_0/dds_state_0/N_534 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[8]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[6]_net_1 ));
    INV \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3_I_4  (
        .A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[0] ));
    AND3 \scalestate_0/necount_cmp_1/AND3_0  (.A(
        \scalestate_0/necount_cmp_1/AND3_1_Y ), .B(
        \scalestate_0/necount_cmp_1/XNOR2_6_Y ), .C(
        \scalestate_0/necount_cmp_1/XNOR2_4_Y ), .Y(
        \scalestate_0/necount_cmp_1/AND3_0_Y ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO_5[3]  (.A(
        \PLUSE_0/bri_state_0/cs[3]_net_1 ), .B(
        \PLUSE_0/bri_state_0/csse_2_0_a4_1_0 ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_0 ));
    MX2B \topctrlchange_0/sw_acq2_RNO_0  (.A(sw_acq2_c), .B(
        \topctrlchange_0/sw_acq2_6_iv ), .S(
        \dds_change_0.un1_change_2 ), .Y(\topctrlchange_0/N_9 ));
    AND2 AND2_0 (.A(Signal_Noise_Acq_0_acq_clk), .B(
        top_code_0_acqclken), .Y(Acq_clk_c));
    NOR2 \scanstate_0/CS_RNIFF4H[6]  (.A(\scanstate_0/CS[7]_net_1 ), 
        .B(\scanstate_0/CS[6]_net_1 ), .Y(\scanstate_0/N_255 ));
    XNOR2 \PLUSE_0/bri_coder_0/half_0_I_1  (.A(\PLUSE_0/half_para[7] ), 
        .B(\PLUSE_0/count_2[7] ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1 \top_code_0/dumpdata[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[3] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_52_i ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_37_i ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_1  (.A(
        \scalestate_0/necount_cmp_0/NOR3A_1_Y ), .B(
        \scalestate_0/necount_cmp_0/OR2A_3_Y ), .C(
        \scalestate_0/necount_cmp_0/NAND3A_3_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_1_Y ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[1]  (.A(
        \ClockManagement_0/long_timer_0/count[1]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[0]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[3]  (
        .D(\s_acq_change_0_s_acqnum[3] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[3]_net_1 )
        );
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_10_RNO_0  
        (.A(\s_acq_change_0_s_stripnum[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N168 ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_10_0 )
        );
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m260  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_261 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m252  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_251 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_252 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_253 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[2]_net_1 ));
    NOR2 \DDS_0/dds_state_0/para_9_i_0_a2_5_0[22]  (.A(\DDS_0/i[0] ), 
        .B(top_code_0_dds_load), .Y(\DDS_0/dds_state_0/N_535_0 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m75  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_76 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[6] ));
    DFN1E1 \scalestate_0/CUTTIME90[19]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[19]_net_1 ));
    DFN1 \DUMP_0/dump_timer_0/count[2]  (.D(
        \DUMP_0/dump_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_1[2] ));
    DFN1E1 \scalestate_0/PLUSETIME180[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[7]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO[16]  (.A(\state_1ms_0/N_83 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[16]_net_1 ));
    NOR3C \scalestate_0/CUTTIME180_448_e  (.A(\scalestate_0/N_60 ), .B(
        \scalestate_0/N_66 ), .C(\top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/N_1661 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[5]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[5] ));
    MX2 \scalestate_0/strippluse_RNO_0[8]  (.A(
        \scalestate_0/strippluse_6[8] ), .B(
        \scalestate_0_strippluse[8] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_567 ));
    OR2 \top_code_0/n_s_ctrl_3_i_o3  (.A(\top_code_0/N_190 ), .B(
        \top_code_0/N_171 ), .Y(\top_code_0/N_198 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_36  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .C(
        \timer_top_0/timer_0/timedata[12]_net_1 ), .Y(
        \timer_top_0/timer_0/N_10 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m163  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_164 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[8]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n8 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_24  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[3] ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[4] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI9O6T[16]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[16]_net_1 ), .B(
        \sd_acq_top_0/count[16] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_16[0] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_25[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[1]_net_1 ), .B(
        \sd_acq_top_0/count_10[1] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_1[0] ));
    OA1 \scalestate_0/timecount_ret_10_RNO  (.A(
        \scalestate_0/N_1153_1 ), .B(\scalestate_0/N_508_i_0_0 ), .C(
        top_code_0_scale_rst_0), .Y(
        \scalestate_0/timecount_cnst_m_0[7] ));
    DFN1E1 \top_code_0/dumpdata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[5] ));
    DFN1E1 \scalestate_0/PLUSETIME90[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[1]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m70_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[0] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI6TN13[14]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_18[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_16[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_3[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_12[0] ));
    DFN1E1 \scalestate_0/CUTTIME180[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[14]_net_1 )
        );
    NOR3C \timer_top_0/timer_0/timedata_RNO[10]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_28_0 ), .Y(
        \timer_top_0/timer_0/timedata_4[10] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m274  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_273 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_274 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_275 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i4_mux ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m45 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_25  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_25_Y ));
    IOPAD_TRI \ddswclk_pad/U0/U0  (.D(\ddswclk_pad/U0/NET1 ), .E(
        \ddswclk_pad/U0/NET2 ), .PAD(ddswclk));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_29  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_29_Y ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[5]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[5] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_1[5] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m44_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[15] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_31  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/timedata[9]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .Y(
        \timer_top_0/timer_0/N_12 ));
    DFN1E1 \scalestate_0/CUTTIME90[4]  (.D(\top_code_0_scaledatain[4] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[4]_net_1 ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_2  (.A(
        \timer_top_0/dataout[2] ), .B(
        \timer_top_0/timer_0/timedata[2]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_2_Y ));
    IOPAD_TRI \relay_on_pad[0]/U0/U0  (.D(\relay_on_pad[0]/U0/NET1 ), 
        .E(\relay_on_pad[0]/U0/NET2 ), .PAD(relay_on[0]));
    DFN1 \PLUSE_0/qq_state_0/cs[4]  (.D(
        \PLUSE_0/qq_state_0/cs_RNO_2[4] ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_0/cs[4]_net_1 ));
    NOR2B \DUMP_ON_0/off_on_timer_0/count_RNIVAKK[2]  (.A(
        \DUMP_ON_0/off_on_timer_0/count_c1 ), .B(
        \DUMP_ON_0/count_5[2] ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_c2 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[19]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[19]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m45_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[14] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[5]  (.D(
        \top_code_0_bri_datain[9] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[5] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[10] ));
    DFN1E1 \noisestate_0/timecount_1[1]  (.D(
        \noisestate_0/timecount_5[1] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m249  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_242 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_249 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[7] ));
    DFN1E1 \top_code_0/pd_pluse_data[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[12] ));
    MX2 \PLUSE_0/bri_timer_0/count[5]/U0  (.A(\PLUSE_0/count_2[5] ), 
        .B(\PLUSE_0/bri_timer_0/count_n5 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[5]/Y ));
    AOI1B \DUMP_OFF_0/off_on_state_0/state_over_RNO_0  (.A(
        \DUMP_OFF_0/off_on_state_0/N_42_i ), .B(
        \DUMP_OFF_0/off_on_state_0_state_over ), .C(
        \DUMP_OFF_0/i_3[0] ), .Y(\DUMP_OFF_0/off_on_state_0/N_12_mux ));
    NOR3A \DUMP_0/dump_state_0/cs_RNO[4]  (.A(
        \DUMP_0/dump_state_0/cs4 ), .B(\DUMP_0/dump_state_0/N_185 ), 
        .C(\DUMP_0/dump_state_0/N_186 ), .Y(
        \DUMP_0/dump_state_0/cs_RNO_0[4]_net_1 ));
    IOPAD_BI \xd_pad[2]/U0/U0  (.D(\xd_pad[2]/U0/NET1 ), .E(
        \xd_pad[2]/U0/NET2 ), .Y(\xd_pad[2]/U0/NET3 ), .PAD(xd[2]));
    DFN1E1 \top_code_0/dds_configdata[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[12] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO[21]  (.A(
        \scalestate_0_timecount[21] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[21]_net_1 ));
    DFN1 \DUMP_0/dump_timer_0/count[3]  (.D(
        \DUMP_0/dump_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_1[3] ));
    OR3 \scalestate_0/timecount_ret_11_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[7] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[7] ), .C(
        \scalestate_0/timecount_20_iv_2[7] ), .Y(
        \scalestate_0/timecount_20_iv_7[7] ));
    DFN1 \scalestate_0/CS[13]  (.D(\scalestate_0/CS_RNO[13]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[13]_net_1 ));
    MX2 \plusestate_0/timecount_1_RNO_0[12]  (.A(
        \plusestate_0/DUMPTIME[12]_net_1 ), .B(
        \plusestate_0/PLUSETIME[12]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_83 ));
    DFN1E1 \bridge_div_0/dataall[0]  (.D(
        \bridge_div_0/DWACT_ADD_CI_0_partial_sum[0] ), .CLK(GLA_net_1), 
        .E(top_code_0_bridge_load), .Q(\bridge_div_0/dataall[0]_net_1 )
        );
    AO1A \scalestate_0/timecount_ret_38_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[3]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[3] ), .Y(
        \scalestate_0/timecount_20_iv_0[3] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m40  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_41_i ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m106  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_107 ));
    NOR2A \DSTimer_0/dump_sustain_timer_0/count_RNO[0]  (.A(
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_n0 ));
    DFN1 \timer_top_0/state_switch_0/dataout[2]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[2]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[2] ));
    XOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIKL7R[3]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[3]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_3 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[11]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c9 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n11 ));
    DFN1E1 \top_code_0/plusedata[13]  (.D(\GPMI_0_dataout[13] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[13] ));
    NOR2B \DDS_0/dds_state_0/para_RNO_1[7]  (.A(
        \DDS_0/dds_state_0/para_reg[7]_net_1 ), .B(
        \DDS_0/dds_state_0/N_535 ), .Y(\DDS_0/dds_state_0/N_272 ));
    AX1C \bridge_div_0/count_5_I_7  (.A(
        \bridge_div_0/count_RNIFNOM7[1]_net_1 ), .B(
        \bridge_div_0/count_RNIEMOM7[0]_net_1 ), .C(
        \bridge_div_0/count_RNIGOOM7[2]_net_1 ), .Y(
        \bridge_div_0/count_5[2] ));
    DFN1E1 \noisestate_0/acqtime[3]  (.D(\top_code_0_noisedata[3] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[3]_net_1 ));
    NOR3B \DUMP_OFF_0/off_on_state_0/cs_RNO[1]  (.A(
        bri_dump_sw_0_reset_out_0), .B(\DUMP_OFF_0/i_3[0] ), .C(
        \DUMP_OFF_0/off_on_state_0/N_10 ), .Y(
        \DUMP_OFF_0/off_on_state_0/cs_nsss[1] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[8]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[8] ));
    OR3 \scalestate_0/timecount_ret_28_RNO_2  (.A(
        \scalestate_0/OPENTIME_m[1] ), .B(
        \scalestate_0/CUTTIME180_m[1] ), .C(
        \scalestate_0/timecount_20_iv_3[1] ), .Y(
        \scalestate_0/timecount_20_iv_7[1] ));
    NOR3A \scalestate_0/CS_RNI73D41[18]  (.A(
        \scalestate_0/un1_CS6_39_i_a2_0 ), .B(\scalestate_0/N_1212 ), 
        .C(\scalestate_0/N_1194 ), .Y(\scalestate_0/N_1304 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m43  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_44 ));
    XOR2 \PLUSE_0/qq_coder_1/i_reg10_0[0]  (.A(\PLUSE_0/qq_para3[0] ), 
        .B(\PLUSE_0/count_7[0] ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_0[0]_net_1 ));
    OA1B \plusestate_0/CS_RNO[3]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[3]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[3] )
        , .Y(\plusestate_0/CS_RNO_0[3]_net_1 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[5]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[5] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[5]_net_1 ));
    OA1B \state_1ms_0/CS_RNO[3]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS[3]_net_1 ), .C(\state_1ms_0/CS_srsts_i_0[3] ), 
        .Y(\state_1ms_0/CS_RNO_3[3] ));
    DFN1E1 \top_code_0/change_0[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/change_1_sqmuxa ), .Q(
        \top_code_0_change_0[1] ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_9  (.A(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .B(
        \timer_top_0/dataout[4] ), .C(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_9_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[0]_net_1 ));
    OR2A \DDS_0/dds_state_0/cs_RNI4SGF_0[6]  (.A(
        \DDS_0/dds_state_0/cs[6]_net_1 ), .B(\DDS_0/i[3] ), .Y(
        \DDS_0/dds_state_0/N_224 ));
    NOR2A \scalestate_0/timecount_RNO_4[20]  (.A(
        \scalestate_0/CUTTIME90[20]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[20] ));
    DFN1E1 \top_code_0/bri_datain[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[11] ));
    NOR3C \scalestate_0/timecount_ret_34_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[9]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[9] ));
    NOR3C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_15[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_i[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[4]_net_1 ));
    AO1A \scalestate_0/timecount_ret_37_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/S_DUMPTIME[3]_net_1 ), .C(
        \scalestate_0/timecount_20_iv_1[3] ), .Y(
        \scalestate_0/timecount_20_iv_6[3] ));
    AO1 \topctrlchange_0/rt_sw_RNO_1  (.A(scalestate_0_rt_sw), .B(
        \top_code_0_change_0[0] ), .C(\topctrlchange_0/rt_swin1_m ), 
        .Y(\topctrlchange_0/rt_sw_6 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m307  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_306 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_307 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_308 ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[5]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_1[5] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[2]  (.A(
        \timer_top_0/state_switch_0/N_232 ), .B(
        \timer_top_0/state_switch_0/N_234 ), .C(
        \timer_top_0/state_switch_0/N_233 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[2] ));
    NOR3C \scalestate_0/timecount_ret_29_RNO_3  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[1]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[1] ));
    DFN1E1 \plusestate_0/DUMPTIME[12]  (.D(\top_code_0_plusedata[12] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[12]_net_1 ));
    MX2 \bri_dump_sw_0/dump_start_RNO_0  (.A(plusestate_0_soft_d), .B(
        scalestate_0_dump_start), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/dump_start_5 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIFAIO1[5]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c4 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c6 ));
    NOR2A \scalestate_0/timecount_ret_20_RNO_4  (.A(
        \scalestate_0/CUTTIME90[8]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[8] ));
    DFN1E1 \top_code_0/state_1ms_lc[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/state_1ms_lc_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_lc[1] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[0]  (.D(
        \top_code_0_sd_sacq_data[0] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[0]_net_1 ));
    DFN1 \DUMP_OFF_0/off_on_state_0/state_over  (.D(
        \DUMP_OFF_0/off_on_state_0/N_9 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/off_on_state_0_state_over ));
    DFN1E1 \top_code_0/state_1ms_data[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[11] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[10]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[10] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_50_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_13[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[2]_net_1 ), .B(
        \sd_acq_top_0/count_10[2] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_2[0] ));
    MX2 \scalestate_0/strippluse_RNO_2[10]  (.A(
        \scalestate_0/STRIPNUM180_NUM[10]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[10]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_430 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[10]  (.A(
        \top_code_0_dumpdata_0[10] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[10] ));
    DFN1E1 \top_code_0/s_acqnum[13]  (.D(\GPMI_0_dataout[13] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[13] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIRG8D[13]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[13]_net_1 )
        , .B(\pd_pluse_top_0/count[13] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_13[0] ));
    NOR2B \top_code_0/relay_on_RNO[0]  (.A(\top_code_0/N_809 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[0]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[7]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[7]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[7]_net_1 )
        );
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI0PEH[15]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[15]_net_1 )
        , .B(\pd_pluse_top_0/count[15] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_15[0] ));
    DFN1 \timer_top_0/state_switch_0/dataout[16]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[16]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[16] ));
    IOPAD_TRI \relay_close_pad[8]/U0/U0  (.D(
        \relay_close_pad[8]/U0/NET1 ), .E(\relay_close_pad[8]/U0/NET2 )
        , .PAD(relay_close[8]));
    XA1C \ClockManagement_0/long_timer_0/timeup_RNO_7  (.A(
        \ClockManagement_0/long_timer_0/count[10]_net_1 ), .B(
        \top_code_0_sigtimedata[10] ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_3 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_6 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_19[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[17]_net_1 ), .B(
        \sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_17[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[10]  (.A(
        \noisestate_0_timecount[10] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_250 ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[9]  (.A(
        \DUMP_0/dump_timer_0/count_c8 ), .B(\DUMP_0/count[9] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n9 ));
    OR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_44_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[1] )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i8_mux ));
    DFN1 \PLUSE_0/qq_state_1/cs[3]  (.D(
        \PLUSE_0/qq_state_1/cs_RNO_2[3] ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_1/cs[3]_net_1 ));
    OA1C \top_code_0/sigrst_RNO  (.A(\top_code_0/N_209 ), .B(
        top_code_0_sigrst), .C(\top_code_0/N_312 ), .Y(
        \top_code_0/N_104 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i18_mux ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIP0JI[8]  (.A(
        \DUMP_0/dump_coder_0/para4[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_8[0] ));
    IOIN_IB \xa_pad[7]/U0/U1  (.YIN(\xa_pad[7]/U0/NET1 ), .Y(\xa_c[7] )
        );
    OA1B \top_code_0/pluse_noise_ctrl_RNO  (.A(\top_code_0/N_147 ), .B(
        \top_code_0/N_176 ), .C(\top_code_0/N_293 ), .Y(
        \top_code_0/N_86 ));
    OR3 \state_1ms_0/timecount_RNO_1[9]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[9] ), .B(
        \state_1ms_0/CUTTIME_m[9] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[9] ), .Y(
        \state_1ms_0/timecount_8[9] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[12]  (.D(
        \top_code_0_state_1ms_data[12] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[12]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_6  (.A(\ADC_c[4] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_1_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_1_net ));
    NOR2B \scalestate_0/strippluse_RNO[7]  (.A(\scalestate_0/N_566 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[7]_net_1 ));
    NOR2A \DDS_0/dds_timer_0/count_RNO[0]  (.A(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .B(\DDS_0/count[0] )
        , .Y(\DDS_0/dds_timer_0/count_n0 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_136  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_160_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_106_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_136_Y ));
    DFN1E1 \top_code_0/n_divnum[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[5] ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_37  (.A(
        \timer_top_0/timer_0/N_10 ), .B(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .Y(
        \timer_top_0/timer_0/I_37_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_13_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_13_net ));
    NOR2B \scalestate_0/strippluse_RNO[8]  (.A(\scalestate_0/N_567 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[8]_net_1 ));
    MX2 \PLUSE_0/bri_timer_0/count[2]/U0  (.A(\PLUSE_0/count_8[2] ), 
        .B(\PLUSE_0/bri_timer_0/count_n2 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[2]/Y ));
    NOR2B \scalestate_0/timecount_ret_57_RNO_0  (.A(
        \scalestate_0/CUTTIME180[0]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[0] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m41_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_ADD_5x5_medium_area_I13_Y  
        (.A(\top_code_0_n_divnum_0[4] ), .B(\top_code_0_n_divnum_0[9] )
        , .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i6_mux ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[4] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[21]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[21]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[0]  (.D(
        \top_code_0_pd_pluse_data[0] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[0]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m273  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_274 ));
    XOR2 \PLUSE_0/qq_coder_1/i_reg10_3[0]  (.A(\PLUSE_0/qq_para3[3] ), 
        .B(\PLUSE_0/count_7[3] ), .Y(
        \PLUSE_0/qq_coder_1/i_reg10_3[0]_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[6]  (
        .D(\s_acq_change_0_s_acqnum[6] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[6]_net_1 )
        );
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[4]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_5[4] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[4]_net_1 ));
    NOR3B \DUMP_OFF_0/off_on_coder_0/i_RNO_0[1]  (.A(
        \DUMP_OFF_0/count_3[4] ), .B(\DUMP_OFF_0/count_3[2] ), .C(
        \DUMP_OFF_0/count_3[3] ), .Y(
        \DUMP_OFF_0/off_on_coder_0/i_0_2[1] ));
    DFN1 \PLUSE_0/qq_coder_0/i[3]  (.D(\PLUSE_0/qq_coder_0/i_RNO_2[3] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_4[3] ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m70  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m70_2 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[10]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[10] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[3] ));
    DFN1 \ClockManagement_0/clk_div500_0/count[3]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[3] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[3]_net_1 ));
    AND3 \scalestate_0/necount_inc_0/AND2_3_inst  (.A(
        \scalestate_0/necount[0]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .C(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/inc_2_net ));
    MX2 \noisestate_0/timecount_1_RNO_0[1]  (.A(
        \noisestate_0/acqtime[1]_net_1 ), .B(
        \noisestate_0/dectime[1]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_58 ));
    DFN1 \s_acq_change_0/s_stripnum[2]  (.D(
        \s_acq_change_0/s_stripnum_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[2] ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_18  (.A(
        \top_code_0_sigtimedata[1] ), .B(
        \ClockManagement_0/long_timer_0/count[1]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_1 ));
    DFN1 \top_code_0/relay_close[7]  (.D(
        \top_code_0/relay_close_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[7] ));
    OR2B \scalestate_0/CS_RNIM5B6[14]  (.A(\scalestate_0/CS[14]_net_1 )
        , .B(top_code_0_scale_rst_4), .Y(\scalestate_0/N_1065 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m81  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_78 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_81 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_82 ));
    MX2 \plusestate_0/timecount_1_RNO_0[13]  (.A(
        \plusestate_0/PLUSETIME[13]_net_1 ), .B(
        \plusestate_0/DUMPTIME[13]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_84 ));
    MX2 \top_code_0/relay_close_RNO_0[7]  (.A(\relay_close_c[7] ), .B(
        \GPMI_0_dataout[7] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_826 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[15]  (.D(
        \top_code_0_state_1ms_data[15] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[15]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m186  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_187 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[0]  (.D(
        \top_code_0_n_acqnum_2[0] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[0]_net_1 ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_13  (.A(
        \scalestate_0/NE_NUM[2]_net_1 ), .B(
        \scalestate_0/necount[2]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_2 ));
    XOR2 \PLUSE_0/qq_coder_0/i_reg10_0[0]  (.A(\PLUSE_0/qq_para3[0] ), 
        .B(\PLUSE_0/count_9[0] ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_0[0]_net_1 ));
    XA1 \DSTimer_0/dump_sustain_timer_0/count_RNO[1]  (.A(
        \DSTimer_0/dump_sustain_timer_0/count[1]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[0]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_n1 ));
    OR2B \top_code_0/un1_state_1ms_rst_n117_18_i_o2_0  (.A(\xa_c[7] ), 
        .B(\xa_c[5] ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_18_i_o2_0_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[5]_net_1 ));
    MX2 \s_acq_change_0/s_rst_RNO_1  (.A(net_33_0), .B(net_45), .S(
        \top_code_0_change_0[0] ), .Y(\s_acq_change_0/s_rst_5 ));
    NOR2B \scalestate_0/necount_RNO[2]  (.A(\scalestate_0/N_732 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[2]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[14]  (.D(
        \top_code_0_pd_pluse_data[14] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[14]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i4_mux ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[12]  (.A(\s_acq_change_0/N_82 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[12]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[7] ));
    DFN1E1 \state_1ms_0/CUTTIME[9]  (.D(\top_code_0_state_1ms_data[9] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[9]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[1]  (.A(
        \top_code_0_dumpdata_0[1] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[1]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_data[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[4] ));
    NOR3A \top_code_0/RAM_Rd_rst_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_164 ), .Y(
        \top_code_0/N_266 ));
    DFN0P0 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[0] ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add )
        , .PRE(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ));
    OR2B \DUMP_0/off_on_state_1/state_over_RNO  (.A(
        \DUMP_0/off_on_state_1/N_12_mux ), .B(
        state1ms_choice_0_reset_out), .Y(\DUMP_0/off_on_state_1/N_9 ));
    DFN1E1 \top_code_0/scalechoice[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0[2] ));
    NOR2B \state_1ms_0/timecount_RNO[2]  (.A(\state_1ms_0/N_69 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[2]_net_1 ));
    AND2 \ClockManagement_0/clk_10k_0/un1_count_1_I_52  (.A(
        \ClockManagement_0/clk_10k_0/count[6]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_pog_array_1_2[0] ));
    NOR3C \PLUSE_0/bri_state_0/cs_RNO_0[3]  (.A(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_6 ), .B(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_5 ), .C(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_10 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_11 ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[4]  (.A(
        \PLUSE_0/bri_state_0/cs[4]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs[3]_net_1 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_RNO_4[4] ));
    NOR3C \scalestate_0/timecount_ret_65_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[13]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[13] ));
    DFN1 \CAL_0/cal_div_0/count[0]  (.D(\CAL_0/cal_div_0/count_5[0] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[0]_net_1 ));
    IOIN_IB \ADC_pad[2]/U0/U1  (.YIN(\ADC_pad[2]/U0/NET1 ), .Y(
        \ADC_c[2] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[11]  (.A(
        \state_1ms_0_timecount[11] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_197 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[2]  (
        .D(\top_code_0_s_periodnum[2] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[2]_net_1 )
        );
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[0]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_9[0] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_10[0] ));
    AO1A \sd_acq_top_0/sd_sacq_state_0/cs_RNIBEGD[12]  (.A(
        \sd_acq_top_0/i[10] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[13]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_230 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_201 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_27  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[2] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[3] )
        );
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[2]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[2] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_5[2] ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_21  (.A(\PLUSE_0/half_para[4] ), 
        .B(\PLUSE_0/count_8[4] ), .Y(\PLUSE_0/bri_coder_0/N_9 ));
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_0  (.A(
        \scalestate_0/necount_cmp_1/NOR3A_0_Y ), .B(
        \scalestate_0/necount_cmp_1/OR2A_5_Y ), .C(
        \scalestate_0/necount_cmp_1/NAND3A_2_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_0_Y ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIGC141[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_22[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_15[0] ));
    DFN1 \DUMP_0/dump_state_0/timer_start  (.D(
        \DUMP_0/dump_state_0/timer_start_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(\DUMP_0/dump_state_0_timer_start ));
    AO1C \DUMP_0/dump_coder_0/un1_para114_3  (.A(
        \DUMP_0/dump_coder_0/para18_net_1 ), .B(
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ), .C(
        top_code_0_dumpload), .Y(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ));
    OR2B \DUMP_0/dump_coder_0/un1_dump_choice_2  (.A(
        \top_code_0_dump_cho_0[2] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ));
    OR2A \PLUSE_0/qq_state_1/cs_RNO_0[1]  (.A(
        \PLUSE_0/qq_state_1/cs[1]_net_1 ), .B(\PLUSE_0/i_7[1] ), .Y(
        \PLUSE_0/qq_state_1/N_82 ));
    MX2 \plusestate_0/timecount_1_RNO_0[5]  (.A(
        \plusestate_0/PLUSETIME[5]_net_1 ), .B(
        \plusestate_0/DUMPTIME[5]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_76 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_30  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[2] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[6] )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m70_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[0] ));
    DFN1P0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/en  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/en_RNO_0 ), 
        .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .PRE(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0_en ));
    OR3 \scalestate_0/timecount_ret_63_RNO  (.A(
        \scalestate_0/CUTTIME180_m[13] ), .B(
        \scalestate_0/OPENTIME_m[13] ), .C(
        \scalestate_0/timecount_20_iv_3[13] ), .Y(
        \scalestate_0/timecount_20_iv_7[13] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m45  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_44 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_45 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_46 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[27]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[27]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_474 ));
    NOR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[2]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_214 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_215 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[2] ));
    NOR3A \dds_change_0/dds_rst_RNO_4  (.A(net_33), .B(
        \top_code_0_change[0] ), .C(\top_code_0_change[1] ), .Y(
        \dds_change_0/ddsrstin1_m ));
    DFN1E1 \plusestate_0/timecount_1[0]  (.D(
        \plusestate_0/timecount_5[0] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[0] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[2]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[2] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIBQ6T[17]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[17]_net_1 ), .B(
        \sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_17[0] ));
    NOR3A \ClockManagement_0/clk_div500_0/count_RNIEA8E1[0]  (.A(
        \ClockManagement_0/clk_5M_en ), .B(
        \ClockManagement_0/clk_div500_0/count[1]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count[0]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_6 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[7]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[8]  (.D(
        \top_code_0_pd_pluse_data[8] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[8]_net_1 ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[4]  (.A(
        \DUMP_0/dump_timer_0/count_c3 ), .B(\DUMP_0/count_1[4] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n4 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[8]  (.D(
        \DUMP_0/dump_coder_0/para2_4[8]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[8]_net_1 ));
    DFN0C0 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[1] ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add )
        , .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[1] ));
    DFN1 \DDS_0/dds_timer_0/count[7]  (.D(\DDS_0/dds_timer_0/count_n7 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[7] ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_1_RNO  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N146 ), 
        .B(\s_acq_change_0_s_stripnum[4] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_4 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[14]  (.D(
        \top_code_0_pd_pluse_data[14] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[14]_net_1 ));
    DFN1E1 \bri_dump_sw_0/turn_delay  (.D(\bri_dump_sw_0/turn_delay_4 )
        , .CLK(GLA_net_1), .E(net_27), .Q(bri_dump_sw_0_turn_delay));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m244  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_243 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_244 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_245 ));
    IOPAD_TRI \cal_out_pad/U0/U0  (.D(\cal_out_pad/U0/NET1 ), .E(
        \cal_out_pad/U0/NET2 ), .PAD(cal_out));
    MX2 \scalestate_0/strippluse_RNO_2[4]  (.A(
        \scalestate_0/STRIPNUM180_NUM[4]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[4]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_424 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_0  (.A(\xd_in[14] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[14] ));
    XO1 \PLUSE_0/qq_coder_0/un1_qq_para2_NE_2[0]  (.A(
        \PLUSE_0/count_9[1] ), .B(\PLUSE_0/qq_para2[1] ), .C(
        \PLUSE_0/qq_coder_0/un1_qq_para2_0[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_NE_2[0]_net_1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_2_RNO_2  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N142 ), 
        .B(\s_acq_change_0_s_stripnum[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_2_0_0 )
        );
    NOR3B \scalestate_0/CUTTIME180_Tini_516_e  (.A(\scalestate_0/N_66 )
        , .B(\scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 ), .C(
        \top_code_0_scalechoice_0_0[0] ), .Y(\scalestate_0/N_1729 ));
    DFN1E1 \scalestate_0/CUTTIME90[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[13]_net_1 ));
    DFN1 \scanstate_0/soft_d  (.D(\scanstate_0/soft_d_RNO_3 ), .CLK(
        GLA_net_1), .Q(scanstate_0_soft_d));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[8] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m226  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_223 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_226 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_227 ));
    AOI1B \DUMP_OFF_1/off_on_state_0/state_over_RNO_0  (.A(
        \DUMP_OFF_1/off_on_state_0/N_42_i ), .B(
        \DUMP_OFF_1/off_on_state_0_state_over ), .C(
        \DUMP_OFF_1/i_4[0] ), .Y(\DUMP_OFF_1/off_on_state_0/N_12_mux ));
    NOR3C \scalestate_0/NE_NUM_1_sqmuxa_0_a2  (.A(
        \top_code_0_scalechoice_0[0] ), .B(\scalestate_0/N_60 ), .C(
        \scalestate_0/N_65 ), .Y(\scalestate_0/NE_NUM_1_sqmuxa ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[8]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_38 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[8] ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m46_3 ));
    XA1C \ClockManagement_0/long_timer_0/timeup_RNO_17  (.A(
        \ClockManagement_0/long_timer_0/count[0]_net_1 ), .B(
        \top_code_0_sigtimedata[0] ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_6 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_4 ));
    DFN1 \timer_top_0/timer_0/timedata[7]  (.D(
        \timer_top_0/timer_0/timedata_4[7] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[7]_net_1 ));
    OR3 \scalestate_0/timecount_ret_59_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[0] ), .B(
        \scalestate_0/OPENTIME_TEL_m[0] ), .C(
        \scalestate_0/timecount_20_iv_4[0] ), .Y(
        \scalestate_0/timecount_20_iv_8[0] ));
    DFN1E1 \scalestate_0/M_NUM[7]  (.D(\top_code_0_scaledatain[7] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[7]_net_1 ));
    NOR3C \PLUSE_0/qq_coder_0/i_RNO_0[1]  (.A(
        bri_dump_sw_0_reset_out_0), .B(\PLUSE_0/qq_coder_0/i_0_1[1] ), 
        .C(\PLUSE_0/qq_coder_0/i_0_2[1] ), .Y(
        \PLUSE_0/qq_coder_0/i_0_4[1] ));
    CLKIO \ddsclkout_pad/U0/U1  (.A(\ddsclkout_pad/U0/NET1 ), .Y(
        ddsclkout_c));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI4PL3E[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_19[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_18[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_127  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_127_Y ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[2]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[2] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[2] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[4]  (.D(
        \top_code_0_state_1ms_data[4] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[4]_net_1 ));
    IOIN_IB \xa_pad[1]/U0/U1  (.YIN(\xa_pad[1]/U0/NET1 ), .Y(\xa_c[1] )
        );
    XOR2 \DUMP_0/dump_coder_0/para6_RNIR6PK[8]  (.A(
        \DUMP_0/dump_coder_0/para6[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_8[0] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m43_1 ));
    OA1C \top_code_0/RAM_Rd_rst_RNO  (.A(\top_code_0/N_206 ), .B(
        top_code_0_RAM_Rd_rst), .C(\top_code_0/N_266 ), .Y(
        \top_code_0/N_58 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m43_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[16] ));
    NOR2B \scalestate_0/strippluse_RNO[2]  (.A(\scalestate_0/N_561 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[2]_net_1 ));
    XA1 \DDS_0/dds_timer_0/count_RNO[3]  (.A(
        \DDS_0/dds_timer_0/count_c2 ), .B(\DDS_0/count[3] ), .C(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DDS_0/dds_timer_0/count_n3 ));
    OR2A \top_code_0/pluse_rst_0_0_RNIO7ND3  (.A(net_27), .B(
        \top_code_0/N_804 ), .Y(
        \top_code_0/pluse_rst_0_0_RNIO7ND3_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I4_un1_CO1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N146 ), 
        .B(\s_acq_change_0_s_stripnum[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I4_un1_CO1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[6] ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI6GTG1[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_26 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_5 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_1 ));
    NOR2B \plusestate_0/dds_config_RNO  (.A(\plusestate_0/N_142 ), .B(
        top_code_0_pluse_rst), .Y(\plusestate_0/dds_config_RNO_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[5]  (.D(
        \DUMP_0/dump_coder_0/para4_4[5]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[5]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_56  (.A(
        \timer_top_0/timer_0/N_4 ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .Y(
        \timer_top_0/timer_0/I_56 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m230  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_231 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/ADD_20x20_slow_I19_Y_4 )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m45 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIQUD42[11]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_14[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_15[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_1[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_8[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m70_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[0] ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_18  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]_net_1 )
        , .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_9 ));
    DFN1E1 \top_code_0/sd_sacq_data[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[2] ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_13  (.A(
        \top_code_0_sigtimedata[5] ), .B(
        \ClockManagement_0/long_timer_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_5 ));
    DFN1 \timer_top_0/timer_0/timedata[3]  (.D(
        \timer_top_0/timer_0/timedata_4[3] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[3]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_51  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[5] ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[28] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m10  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i4_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[3] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i6_mux ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_2  (.A(
        \timer_top_0/dataout[17] ), .B(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_2_Y ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[9] ));
    NOR3A \scalestate_0/intertodsp_RNO_2  (.A(\scalestate_0/N_1269 ), 
        .B(\scalestate_0/CS[16]_net_1 ), .C(\scalestate_0/N_1210 ), .Y(
        \scalestate_0/un1_CS_27 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i4_mux ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_RNO  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop ), .B(
        scan_scale_sw_0_s_start), .C(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_RNO_net_1 )
        );
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_0  (.A(
        \scalestate_0/M_NUM[3]_net_1 ), .B(
        \scalestate_0/necount[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_0_Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m10  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_9_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_10_0 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_11_0 ));
    DFN1 \s_acq_change_0/s_acqnum[11]  (.D(
        \s_acq_change_0/s_acqnum_RNO[11]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[11] ));
    NOR3C \scalestate_0/OPENTIME_468_e  (.A(\scalestate_0/N_62 ), .B(
        \scalestate_0/N_65 ), .C(\top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/N_1681 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m133  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_132 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_133 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_134 ));
    DFN1 \scanstate_0/CS[7]  (.D(\scanstate_0/CS_RNO_2[7] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[7]_net_1 ));
    DFN1 \scalestate_0/CS[17]  (.D(\scalestate_0/CS_RNO[17]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[17]_net_1 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[3]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m128  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[19] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_129 ));
    XO1 \DUMP_0/dump_coder_0/para2_RNIGNP01[9]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_coder_0/para2[9]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_3_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_5[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_8_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_30_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_152_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_8_inst ));
    DFN1E1 \scalestate_0/PLUSETIME90[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[3]_net_1 ));
    DFN1E1 \plusestate_0/DUMPTIME[1]  (.D(\top_code_0_plusedata[1] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[1]_net_1 ));
    DFN1E1 \top_code_0/dumpdata[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[1] ));
    MX2 \scanstate_0/timecount_1_RNO_0[10]  (.A(
        \scanstate_0/acqtime[10]_net_1 ), .B(
        \scanstate_0/dectime[10]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_68 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m105  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_106 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[5] ));
    NOR3B \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[0]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/count_6[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[0] ));
    DFN1E1 \top_code_0/scandata[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[10] ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[6]  (.A(
        \s_acq_change_0/s_stripnum_5[6] ), .B(
        \s_acq_change_0_s_stripnum[6] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_62 ));
    NOR3A \DUMP_0/dump_coder_0/para17  (.A(\top_code_0_dump_cho_0[1] ), 
        .B(\top_code_0_dump_cho_0[2] ), .C(\top_code_0_dump_cho_0[0] ), 
        .Y(\DUMP_0/dump_coder_0/para17_net_1 ));
    MX2 \state1ms_choice_0/reset_out_RNO_0  (.A(
        bri_dump_sw_0_reset_out_0), .B(state_1ms_0_reset_out), .S(
        top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/reset_out_5 ));
    DFN1 \scalestate_0/CS[10]  (.D(\scalestate_0/CS_RNO[10]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[10]_net_1 ));
    IOPAD_TRI \s_acq180_pad/U0/U0  (.D(\s_acq180_pad/U0/NET1 ), .E(
        \s_acq180_pad/U0/NET2 ), .PAD(s_acq180));
    NOR2B \state_1ms_0/soft_dump_RNO  (.A(\state_1ms_0/N_152 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/soft_dump_RNO_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m8  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[17] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_9_0 ));
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_42  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[7] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[8] ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[5] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[10] ));
    MX2 \state_1ms_0/timecount_RNO_0[1]  (.A(
        \state_1ms_0/timecount_8[1] ), .B(\state_1ms_0_timecount[1] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_68 ));
    DFN1E1 \scanstate_0/timecount_1[9]  (.D(
        \scanstate_0/timecount_5[9] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[9] ));
    AO1B \PLUSE_0/qq_state_0/stateover_RNO  (.A(
        \PLUSE_0/qq_state_0_stateover ), .B(\PLUSE_0/qq_state_0/N_84 ), 
        .C(\PLUSE_0/qq_state_0/cs4 ), .Y(
        \PLUSE_0/qq_state_0/stateover_RNO_0 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[15]  (.D(
        \top_code_0_state_1ms_data[15] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[15]_net_1 ));
    OA1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_62  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6_0 ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8_0 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7_0 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_11_0 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i12_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_76  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_101_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_60_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_76_Y ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[8]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c6 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n8 ));
    NOR2B \scalestate_0/timecount_ret_52_RNO  (.A(
        \scalestate_0/OPENTIME_TEL[18]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[18] ));
    XOR2 \bridge_div_0/dataall_RNIA2OO[3]  (.A(
        \bridge_div_0/dataall[3]_net_1 ), .B(
        \bridge_div_0/count[3]_net_1 ), .Y(
        \bridge_div_0/un1_count_3[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_131  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_131_Y ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m243  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_244 ));
    DFN1E1 \scanstate_0/dectime[0]  (.D(\top_code_0_scandata[0] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[0]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[9]  (.D(
        \DUMP_0/dump_coder_0/para4_4[9]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[9]_net_1 ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/data_RNO[0]  (.A(
        \DSTimer_0/dump_sustain_timer_0/N_24 ), .B(
        top_code_0_dump_sustain), .Y(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[0]_net_1 ));
    DFN1 \s_acq_change_0/s_acqnum[14]  (.D(
        \s_acq_change_0/s_acqnum_RNO[14]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[14] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[11]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[11] ));
    NOR3A \topctrlchange_0/soft_dump_6_iv_RNO_1  (.A(
        nsctrl_choice_0_soft_d), .B(\top_code_0_change_0[0] ), .C(
        \top_code_0_change[1] ), .Y(\topctrlchange_0/s_dumpin1_m ));
    DFN1E1 \scalestate_0/timecount_ret_37  (.D(
        \scalestate_0/timecount_20_iv_6[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[3] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[27]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[27]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_475 ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_6  (.A(
        \top_code_0_sigtimedata[7] ), .B(
        \ClockManagement_0/long_timer_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_7 ));
    AND3C \top_code_0/un1_state_1ms_rst_n117_4_i_a2  (.A(
        \top_code_0/N_144 ), .B(\top_code_0/N_161 ), .C(
        \top_code_0/N_171 ), .Y(\top_code_0/N_258 ));
    AO1C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_9  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[3]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_5 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[2]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[2]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_8[2] ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[3]  (.D(
        \DUMP_0/dump_coder_0/para4_4[3]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[3]_net_1 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_52  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[3] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[6] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[10] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] )
        );
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNIFKA5[8]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c6 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c8 ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_12  (.A(
        \timer_top_0/dataout[11] ), .B(
        \timer_top_0/timer_0/timedata[11]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_12_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_41  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_41_Y ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[1]  (.A(
        \scalestate_0/ACQ180_NUM[1]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[1]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_449 ));
    MX2 \scalestate_0/strippluse_RNO_2[7]  (.A(
        \scalestate_0/STRIPNUM180_NUM[7]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[7]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_427 ));
    DFN1C0 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10]/U1  (
        .D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ));
    NOR2A \scalestate_0/CS_RNO[21]  (.A(top_code_0_scale_rst_5), .B(
        \scalestate_0/N_1236 ), .Y(\scalestate_0/CS_RNO[21]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[5]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[5] ));
    NOR2A \DDS_0/dds_state_0/para_reg_69_e  (.A(top_code_0_dds_load), 
        .B(top_code_0_dds_choice), .Y(\DDS_0/dds_state_0/N_538 ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIOTFH[8]  (.A(
        \DUMP_0/dump_coder_0/para3[8]_net_1 ), .B(\DUMP_0/count[8] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_8[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[1]_net_1 ));
    NOR2A \scalestate_0/timecount_ret_91_RNO_1  (.A(
        \scalestate_0/DUMPTIME[8]_net_1 ), .B(\scalestate_0/N_1093 ), 
        .Y(\scalestate_0/DUMPTIME_m[8] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[0]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/un1_noise_addr_1_i[0] )
        , .CLK(\Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i16_mux ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[4]  (.D(
        \ClockManagement_0/long_timer_0/count_n4 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[4]_net_1 ));
    NOR3A \top_code_0/pd_pluse_data_1_sqmuxa_0_a2  (.A(
        \top_code_0/dds_configdata_1_sqmuxa_1 ), .B(\top_code_0/N_150 )
        , .C(\top_code_0/N_167 ), .Y(
        \top_code_0/pd_pluse_data_1_sqmuxa ));
    AND2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_14_inst  
        (.A(\pd_pluse_top_0/count[12] ), .B(\pd_pluse_top_0/count[13] )
        , .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_20_net ));
    DFN1 \CAL_0/cal_div_0/cal  (.D(\CAL_0/cal_div_0/cal_RNO_net_1 ), 
        .CLK(ddsclkout_c), .Q(cal_out_c));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[12]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[12]_net_1 ), .CLK(
        ddsclkout_c), .Q(\sd_acq_top_0/sd_sacq_state_0/cs[12]_net_1 ));
    NOR3C \timer_top_0/state_switch_0/clk_en_scale_0_0_a6_0_a5  (.A(
        net_27), .B(\timer_top_0/timer_0_time_up ), .C(
        top_code_0_scale_start), .Y(
        \timer_top_0/state_switch_0/clk_en_scale_0_0_a6_0_a5_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_5[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[3]_net_1 ), .B(
        \pd_pluse_top_0/count_6[3] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_3[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[2]  (.D(
        \DUMP_0/dump_coder_0/para4_4[2]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[2]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[1]_net_1 ));
    OA1 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_21  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_11 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_10 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[0] )
        );
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_9_inst  
        (.A(\pd_pluse_top_0/count_1[6] ), .B(
        \pd_pluse_top_0/count_1[7] ), .C(\pd_pluse_top_0/count_0[8] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net )
        );
    NOR3A \top_code_0/sigtimedata_1_sqmuxa_0_a2  (.A(
        \top_code_0/sigtimedata_1_sqmuxa_1 ), .B(\top_code_0/N_151 ), 
        .C(\top_code_0/N_158 ), .Y(\top_code_0/sigtimedata_1_sqmuxa ));
    DFN1E1 \top_code_0/dump_sustain_data[0]  (.D(\GPMI_0_dataout[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dump_sustain_data_1_sqmuxa ), 
        .Q(\top_code_0_dump_sustain_data[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[5]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[15]_net_1 ));
    NOR2 \scalestate_0/timecount_ret_7_RNO  (.A(
        \scalestate_0/CS[16]_net_1 ), .B(\scalestate_0/N_1206 ), .Y(
        \scalestate_0/timecount_cnst_m_0[3] ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_57  (.A(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[14] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_54_i ));
    OA1B \top_code_0/pluse_lc_RNO_0  (.A(\top_code_0/N_149 ), .B(
        \top_code_0/N_175 ), .C(top_code_0_pluse_lc), .Y(
        \top_code_0/N_291 ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNIFMII[3]  (.A(
        \DUMP_0/dump_coder_0/para4[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_3[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[17]  (.A(
        \scalestate_0_timecount[17] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_268 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[1]  (.A(
        \Signal_Noise_Acq_0/un1_signal_acq_0[1] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_1_inst ), .S(top_code_0_n_s_ctrl_0), 
        .Y(\Signal_Noise_Acq_0_dataout[1] ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_16  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[1] )
        );
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[1]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m18  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_15_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_18_0 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_19_0 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_37  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_37_Y ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[1]  (.A(\scalestate_0/N_449 ), 
        .B(\scalestate_0/ACQECHO_NUM[1]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[1] ));
    DFN1E1 \scalestate_0/CUTTIME180[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[6]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIL0PK[5]  (.A(
        \DUMP_0/dump_coder_0/para6[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_5[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m269  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_270 ));
    IOBI_IB_OB_EB \xd_pad[2]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[2] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[2]/U0/NET3 ), .DOUT(\xd_pad[2]/U0/NET1 ), .EOUT(
        \xd_pad[2]/U0/NET2 ), .Y(\xd_in[2] ));
    NOR2A \noisestate_0/timecount_1_RNO[10]  (.A(\noisestate_0/N_67 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[10] ));
    DFN1E1 \top_code_0/n_acqnum[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[10] ));
    AO1C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_7  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[2]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_0 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_8 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/HOR2_10_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_13_net ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[13] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m45_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[14] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[9]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[9] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_0[9] ));
    AO1 \state_1ms_0/timecount_RNO_4[0]  (.A(
        \state_1ms_0/S_DUMPTIME[0]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[0] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m91  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[5] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_92 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[21]  (.A(
        \DDS_0/dds_state_0/N_512 ), .B(\DDS_0/dds_state_0/N_511 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[21] ), .Y(
        \DDS_0/dds_state_0/N_167 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m250  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[15] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_251 ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_5  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_8_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_3_Y ), .C(
        \timer_top_0/dataout[12] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_5_Y ));
    NOR2A \timer_top_0/state_switch_0/state_start5_0_0_a2_12  (.A(
        net_27), .B(top_code_0_pluse_str), .Y(
        \timer_top_0/state_switch_0/N_282 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[3]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[3] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_6[3] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_139  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_84_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_46_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_139_Y ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m47_4 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_32  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_162_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_105_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_32_Y ));
    NOR2B \bri_dump_sw_0/pluse_start_RNO  (.A(
        \bri_dump_sw_0/pluse_start_5 ), .B(net_27), .Y(
        \bri_dump_sw_0/pluse_start_RNO_net_1 ));
    AO1B \plusestate_0/state_over_n_RNO  (.A(plusestate_0_state_over_n)
        , .B(\plusestate_0/N_302 ), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/state_over_n_RNO_0 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m185  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_186 ));
    DFN1E1 \scalestate_0/timecount_ret_32  (.D(
        \scalestate_0/timecount_20_iv_8[4]_net_1 ), .CLK(GLA_net_1), 
        .E(\scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[4] ));
    AO1 \PLUSE_0/bri_coder_0/un2lto7_2  (.A(\PLUSE_0/count_8[2] ), .B(
        \PLUSE_0/count_8[1] ), .C(\PLUSE_0/count_8[4] ), .Y(
        \PLUSE_0/bri_coder_0/un2lto7_2_net_1 ));
    XA1 \DUMP_0/off_on_timer_0/count_RNO[3]  (.A(\DUMP_0/count_2[3] ), 
        .B(\DUMP_0/off_on_timer_0/count_c2 ), .C(
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_0/count_n3 ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[8] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_6 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[8]_net_1 ));
    XA1A \scalestate_0/necount_cmp_1/AND2_0  (.A(
        \scalestate_0/NE_NUM[9]_net_1 ), .B(
        \scalestate_0/necount[9]_net_1 ), .C(
        \scalestate_0/necount_cmp_1/XNOR2_1_Y ), .Y(
        \scalestate_0/necount_cmp_1/AND2_0_Y ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[1]  (.A(
        \PLUSE_0/bri_state_0/cs[1]_net_1 ), .B(
        \PLUSE_0/bri_state_0/csse_0_0_0_tz ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[1] ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[10]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[10]_net_1 ), .CLK(
        ddsclkout_c), .Q(
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI0ENS[10]  (.A(
        \sd_acq_top_0/count_1[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[10]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_6[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_5[0] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[3]  (.A(
        \scalestate_0/ACQ180_NUM[3]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[3]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_451 ));
    DFN1E0 \DDS_0/dds_state_0/para[22]  (.D(\DDS_0/dds_state_0/N_40 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[22]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m153  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_152 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_153 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_154 ));
    AO1 \scalestate_0/timecount_ret_48_RNO  (.A(
        \scalestate_0/OPENTIME[17]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[17] ), .Y(
        \scalestate_0/timecount_20_0_iv_0[17] ));
    DFN1E1 \scanstate_0/timecount_1[4]  (.D(
        \scanstate_0/timecount_5[4] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[4] ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_15  (.A(
        \top_code_0_sigtimedata[14] ), .B(
        \ClockManagement_0/long_timer_0/count[14]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_14 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[7]  (.D(
        \top_code_0_state_1ms_data[7] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[7]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[1]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[1] ));
    DFN1E1 \state_1ms_0/PLUSETIME[12]  (.D(
        \top_code_0_state_1ms_data[12] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[12]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_78  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_78_Y ));
    DFN1E1 \top_code_0/n_divnum[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[0] ));
    DFN1 \s_acq_change_0/s_stripnum[8]  (.D(
        \s_acq_change_0/s_stripnum_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[8] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[8]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[8] ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[4]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[4] ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[4]_net_1 )
        );
    OA1B \noisestate_0/CS_RNO[2]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[2]_net_1 ), .C(\noisestate_0/CS_srsts_i_0[2] )
        , .Y(\noisestate_0/CS_RNO[2]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[1]  (.D(\GPMI_0_dataout[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[1] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[9]  (.A(
        \scalestate_0_timecount[9] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_203 ));
    AO1 \state_1ms_0/timecount_RNO_2[11]  (.A(
        \state_1ms_0/M_DUMPTIME[11]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[11] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[11] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNISV421[1]  (.A(
        \sd_acq_top_0/count_10[1] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[1]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_5[0] ));
    NOR2 \PLUSE_0/bri_state_0/cs_RNO_8[3]  (.A(
        \PLUSE_0/bri_state_0/cs[5]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs[9]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_3 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[8]  (.D(\top_code_0_scaledatain[8] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[8]_net_1 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[4]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[4]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_8[4] ));
    NOR3A \state_1ms_0/PLUSECYCLE_0_sqmuxa_0_a2  (.A(
        \state_1ms_0/N_17 ), .B(\top_code_0_state_1ms_lc[0] ), .C(
        \top_code_0_state_1ms_lc[1] ), .Y(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIG8A71[14]  (.A(
        \sd_acq_top_0/count_0[14] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[14]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_8[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_3[0] ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[6]  (.A(\scalestate_0/N_553 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[6]_net_1 ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[11]_net_1 ));
    DFN1 \DUMP_OFF_0/off_on_timer_0/count[0]  (.D(
        \DUMP_OFF_0/off_on_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/count_3[0] ));
    DFN1E1 \scalestate_0/timecount_ret_49  (.D(
        \scalestate_0/OPENTIME_TEL_m[17] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/OPENTIME_TEL_m_reto[17] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_13_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_13_net ));
    IOTRI_ORE_EB \soft_dump_pad/U0/U1  (.D(
        \state1ms_choice_0/soft_dump_4 ), .E(VCC), .OCE(net_27), .OCLK(
        GLA_net_1), .DOUT(\soft_dump_pad/U0/NET1 ), .EOUT(
        \soft_dump_pad/U0/NET2 ));
    DFN1E1 \scalestate_0/OPENTIME[9]  (.D(\top_code_0_scaledatain[9] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[9]_net_1 ));
    DFN1E1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[0]  
        (.D(\top_code_0_s_periodnum[0] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[0]_net_1 )
        );
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m46_6 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i10_mux ));
    OR3 \scalestate_0/timecount_ret_20_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[8] ), .B(
        \scalestate_0/OPENTIME_TEL_m[8] ), .C(
        \scalestate_0/timecount_20_iv_4[8] ), .Y(
        \scalestate_0/timecount_20_iv_8[8] ));
    DFN1E1 \scanstate_0/acqtime[8]  (.D(\top_code_0_scandata[8] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[8]_net_1 ));
    NOR3A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_8[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_3[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_1[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_12[4] ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y ));
    OR3B \DUMP_0/dump_coder_0/un1_para114  (.A(
        \top_code_0_dump_cho_0[2] ), .B(top_code_0_dumpload), .C(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ));
    NOR3C \scalestate_0/timecount_ret_70_RNO_1  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[15]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[15] ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNISEG11[11]  
        (.A(\pd_pluse_top_0/count_0[11] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[11]_net_1 ), 
        .C(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_8[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_1[0] ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_49  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_50_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[7] )
        );
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_RNI2MLE  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_net_1 ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0_Signal_acq_clk ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i8_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[11]_net_1 ));
    DFN1 \scalestate_0/CS[4]  (.D(\scalestate_0/CS_RNO_1[4] ), .CLK(
        GLA_net_1), .Q(\scalestate_0/CS[4]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_104  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_104_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI34N5[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_6[0] ));
    AO1A \scalestate_0/timecount_ret_62_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[12]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[12] ), .Y(
        \scalestate_0/timecount_20_iv_0[12] ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[7]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_36 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[7] ));
    DFN1E1 \scalestate_0/PLUSETIME90[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[12]_net_1 ));
    IOPAD_BI \xd_pad[8]/U0/U0  (.D(\xd_pad[8]/U0/NET1 ), .E(
        \xd_pad[8]/U0/NET2 ), .Y(\xd_pad[8]/U0/NET3 ), .PAD(xd[8]));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i22_mux ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y ));
    NOR3C \scalestate_0/timecount_ret_20_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[8]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[8] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[11]  (.A(
        \top_code_0_s_acqnum_2[11] ), .B(\scalestate_0_s_acqnum[11] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[11] ));
    DFN1 \scalestate_0/CS_i[0]  (.D(\scalestate_0/CS_i_RNO_0[0] ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS_i[0]_net_1 ));
    NOR2B \DUMP_0/dump_coder_0/i_RNO[1]  (.A(bri_div_start_0), .B(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/dump_coder_0/i_RNO_0[1] ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[5]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_32_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[5] ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[3]  (.A(
        \top_code_0_dumpdata_0[3] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[3]_net_1 ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_13  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[7]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_4 ));
    AOI1 \scalestate_0/CS_RNO[8]  (.A(\scalestate_0/N_1209_0 ), .B(
        timer_top_0_clk_en_scale_0), .C(\scalestate_0/CS_srsts_i_0[8] )
        , .Y(\scalestate_0/CS_RNO_0[8]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_62_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[12]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[12] ));
    AND3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_10  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/DWACT_FINC_E[0] )
        );
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[4]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c2 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n4 ));
    NOR3A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_6[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_6[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_11[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_14[10] ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_4_inst  (.A(
        \scalestate_0/necount_inc_0/Rcout_5_net ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount1[5] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[3]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c2 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n3 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m41  
        (.A(\s_acq_change_0_s_stripnum[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[11]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i20_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_42_i ));
    DFN1 \scalestate_0/M_pulse  (.D(\scalestate_0/M_pulse_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/M_pulse_net_1 ));
    NOR3C \ClockManagement_0/clk_div500_0/count_RNIA33G1[5]  (.A(
        \ClockManagement_0/clk_div500_0/count[5]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[4]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_2 ), .Y(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa_5 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[8]  (.D(
        \top_code_0_state_1ms_data[8] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[8]_net_1 ));
    NOR2B \scalestate_0/necount_LE_M_RNIMMTM  (.A(
        \scalestate_0/timecount_12_sqmuxa_0 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/N_258 ));
    DFN1 \ClockManagement_0/long_timer_0/clk_5K_reg2  (.D(
        \ClockManagement_0/long_timer_0/clk_5K_reg2_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(
        \ClockManagement_0/long_timer_0/clk_5K_reg2_net_1 ));
    MX2A \scalestate_0/CS_RNO_0[13]  (.A(\scalestate_0/CS[13]_net_1 ), 
        .B(\scalestate_0/N_1195 ), .S(timer_top_0_clk_en_scale_0), .Y(
        \scalestate_0/N_1237 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m59  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[0] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_60 ));
    AND2 \bridge_div_0/dataall_1_I_5  (.A(\top_code_0_scaleddsdiv[1] ), 
        .B(\top_code_0_scaleddsdiv[4] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_1[0] ));
    IOPAD_TRI \sw_acq1_pad/U0/U0  (.D(\sw_acq1_pad/U0/NET1 ), .E(
        \sw_acq1_pad/U0/NET2 ), .PAD(sw_acq1));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m42_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[17] ));
    OR3 \scalestate_0/timecount_ret_69_RNIJ9I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[15] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[15] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[15] ), .Y(
        \scalestate_0_timecount[15] ));
    NOR3C \scalestate_0/timecount_ret_62_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[12]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[12] ));
    NOR2B \top_code_0/relay_close_RNO[9]  (.A(\top_code_0/N_828 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[9]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_29  (.A(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[5] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[2]  (.D(
        \top_code_0_bri_datain[6] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[2] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_56_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI25Q6[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_5[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m47_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] ));
    DFN1E1 \scalestate_0/timecount_ret_1  (.D(
        \scalestate_0/timecount_20_iv_9[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_9_reto[5] ));
    DFN1E1 \scalestate_0/M_NUM[1]  (.D(\top_code_0_scaledatain_0[1] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[1]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m43_2 ));
    AO1 \scalestate_0/timecount_20_iv_5[4]  (.A(
        \scalestate_0/OPENTIME_TEL[4]_net_1 ), .B(\scalestate_0/N_258 )
        , .C(\scalestate_0/timecount_20_iv_0[4] ), .Y(
        \scalestate_0/timecount_20_iv_5[4]_net_1 ));
    DFN1 \ClockManagement_0/clk_10k_0/count[8]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[8] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[8]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[11]  (.A(
        \state_1ms_0/PLUSECYCLE[11]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[11] ));
    NOR2 \syn_md_module_1/syn_md_combine_0/syn_md_temp_0  (.A(
        scalestate_0_sw_acq2), .B(scalestate_0_soft_d), .Y(
        \syn_md_module_1/syn_md_combine_0/syn_md_temp_0_net_1 ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI7RDFA[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_10 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_9 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_11 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE ));
    DFN1E1 \top_code_0/s_addchoice[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice[3] ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[1]  (.D(
        \top_code_0_state_1ms_data[1] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[1]_net_1 ));
    DFN1E0 \DDS_0/dds_state_0/para[27]  (.D(\DDS_0/dds_state_0/N_127 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[27]_net_1 ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_2  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_9_0 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_3 )
        );
    DFN1E1 \top_code_0/dds_load  (.D(\top_code_0/N_68 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_dds_load));
    NOR2B \s_acq_change_0/s_acqnum_RNO[1]  (.A(\s_acq_change_0/N_71 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[1]_net_1 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[11]  (.A(
        \timer_top_0/state_switch_0/N_195 ), .B(
        \timer_top_0/state_switch_0/N_196 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[11] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[11]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[1]  (.A(
        \top_code_0_dumpdata_0[1] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[1]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[11] ));
    AO1A \scalestate_0/necount_LE_M_RNIB1CB1  (.A(
        \scalestate_0/necount_LE_M_RNIBQQD_net_1 ), .B(
        top_code_0_scale_rst_1), .C(\scalestate_0/N_259 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_7_0 ));
    AND3 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/TAND2_15_inst  
        (.A(\pd_pluse_top_0/count[12] ), .B(\pd_pluse_top_0/count[13] )
        , .C(\pd_pluse_top_0/count[14] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_22_net ));
    NOR2 \PLUSE_0/qq_state_1/cs_RNO_1[2]  (.A(\PLUSE_0/i_7[1] ), .B(
        Q4Q5_c), .Y(\PLUSE_0/qq_state_1/N_88 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[11]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[11] ));
    MX2 \PLUSE_0/bri_coder_0/i[3]/U0  (.A(\PLUSE_0/i_3[3] ), .B(net_51)
        , .S(clk_4f_en_0), .Y(\PLUSE_0/bri_coder_0/i[3]/Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m127  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_120 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_127 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_128 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/VAND2_18_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_24_net ), 
        .C(\sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_16_net ));
    DFN1E1 \scalestate_0/CUTTIME180[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[11]_net_1 )
        );
    NOR2A \DUMP_OFF_1/off_on_timer_0/count_RNO[0]  (.A(
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DUMP_OFF_1/count_4[0] ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_n0 ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/data_RNO[2]  (.A(
        \DSTimer_0/dump_sustain_timer_0/N_26 ), .B(
        top_code_0_dump_sustain), .Y(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[2]_net_1 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_7  (.A(
        \timer_top_0/dataout[18] ), .B(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_7_Y ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[7]  (.A(\s_acq_change_0/N_77 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[7]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[8] ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIFBGQ[8]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_6 ), .B(
        \s_acq_change_0_s_stripnum[8] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[8]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_8 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i16_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[2]_net_1 ));
    NOR2B \scanstate_0/soft_d_RNO  (.A(\scanstate_0/N_110 ), .B(net_33)
        , .Y(\scanstate_0/soft_d_RNO_3 ));
    DFN1E1 \scalestate_0/timecount_ret_73  (.D(
        \scalestate_0/timecount_20_iv_8[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[7] ));
    OA1A \scalestate_0/dumpoff_ctr_RNO  (.A(\scalestate_0/N_1187 ), .B(
        scalestate_0_dumpoff_ctr), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/dumpoff_ctr_RNO_2 ));
    NOR3B \top_code_0/s_acqnum_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/s_acqnum_1_sqmuxa_1 ), .C(\top_code_0/N_152 ), .Y(
        \top_code_0/s_acqnum_1_sqmuxa ));
    NOR3B \scalestate_0/ACQECHO_NUM_1_sqmuxa_0_a2_0  (.A(
        top_code_0_scaleload), .B(\top_code_0_scalechoice_0[1] ), .C(
        \top_code_0_scalechoice_0[4] ), .Y(\scalestate_0/N_60 ));
    DFN1E1 \scalestate_0/timecount_ret_69  (.D(
        \scalestate_0/timecount_20_iv_7[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[15] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m43_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI2E811[15]  (.A(
        \sd_acq_top_0/count_0[15] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[15]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_12[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_4[0] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[2]  (.D(
        \top_code_0_pd_pluse_data[2] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[2]_net_1 ));
    AO1C \scalestate_0/pluse_start_RNO_1  (.A(\scalestate_0/N_1197 ), 
        .B(\scalestate_0/N_1263 ), .C(timer_top_0_clk_en_scale), .Y(
        \scalestate_0/N_1171 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m49  
        (.A(\s_acq_change_0_s_stripnum[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[7]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i12_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_50_i ));
    DFN1E1 \top_code_0/n_divnum[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[6] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[8]  (.A(
        \scalestate_0_timecount[8] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_248 ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa_0_a2_0  
        (.A(\top_code_0_sd_sacq_choice[1] ), .B(
        \top_code_0_sd_sacq_choice[3] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_24 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[5]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[8]  (.A(
        \top_code_0_dumpdata_0[8] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[8]_net_1 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_39  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_54_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[0] )
        );
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m303  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] ), .C(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_304 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m28  
        (.A(\s_acq_change_0_s_stripnum[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[9]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i18_mux )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i20_mux ));
    OR3 \scalestate_0/timecount_ret_5_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[2] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[2] ), .C(
        \scalestate_0/timecount_20_iv_2[2] ), .Y(
        \scalestate_0/timecount_20_iv_7[2] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m9  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[1] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_10_0 ));
    DFN1 \DUMP_OFF_0/off_on_state_0/cs[0]  (.D(
        \DUMP_OFF_0/off_on_state_0/N_36_i ), .CLK(GLA_net_1), .Q(
        DUMP_OFF_0_dump_off));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m264  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_257 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_264 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[15] ));
    MX2 \plusestate_0/timecount_1_RNO_0[2]  (.A(
        \plusestate_0/DUMPTIME[2]_net_1 ), .B(
        \plusestate_0/PLUSETIME[2]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_73 ));
    NOR3A \top_code_0/bridge_load_3_i_a2_0  (.A(\top_code_0/N_333 ), 
        .B(\top_code_0/N_144 ), .C(\top_code_0/N_148 ), .Y(
        \top_code_0/N_270 ));
    NOR2B \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[1]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[8]_net_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[1] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_22  (.A(
        \timer_top_0/dataout[8] ), .B(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_22_Y ));
    NOR2A \plusestate_0/DUMPTIME_0_sqmuxa  (.A(top_code_0_pluseload), 
        .B(top_code_0_pluse_lc), .Y(
        \plusestate_0/DUMPTIME_0_sqmuxa_net_1 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m31  
        (.A(\s_acq_change_0_s_stripnum[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[10]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i20_mux )
        );
    OA1B \top_code_0/pluse_scale_RNO  (.A(\top_code_0/N_157 ), .B(
        \top_code_0/N_176 ), .C(\top_code_0/N_295 ), .Y(
        \top_code_0/N_88 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[21]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_62 ), .Y(
        \timer_top_0/timer_0/timedata_4[21] ));
    DFN1 \state_1ms_0/bri_cycle  (.D(
        \state_1ms_0/bri_cycle_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        state_1ms_0_bri_cycle));
    OAI1 \plusestate_0/CS_RNI1ON21[9]  (.A(\plusestate_0/CS[5]_net_1 ), 
        .B(\plusestate_0/CS[9]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/N_271 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[9] ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[3] ), .CLK(
        GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 ));
    OR3 \PLUSE_0/qq_coder_1/un1_qq_para2_NE[0]  (.A(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_1[0]_net_1 ), .B(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_0[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_1/un1_qq_para2_NE_2[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_i[0] ));
    OR2 \top_code_0/sigtimedata_1_sqmuxa_0_o2_0  (.A(\xa_c[3] ), .B(
        \xa_c[2] ), .Y(\top_code_0/N_158 ));
    DFN1 \plusestate_0/CS[1]  (.D(\plusestate_0/CS_RNO_0[1]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[1]_net_1 ));
    DFN1 \s_acq_change_0/s_load_0_0  (.D(
        \s_acq_change_0/s_load_0_0_RNIEJ0I1_net_1 ), .CLK(GLA_net_1), 
        .Q(s_acq_change_0_s_load_0));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[1] ));
    NOR3B \top_code_0/dumpdata_1_sqmuxa_0_a2  (.A(\top_code_0/N_331 ), 
        .B(\top_code_0/N_334 ), .C(\top_code_0/N_159 ), .Y(
        \top_code_0/dumpdata_1_sqmuxa ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[10]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[10] ));
    XO1 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNI25FM1[2]  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[2]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_1 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE_1 ));
    XO1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI5TMK[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_60_i ));
    NOR2B \scalestate_0/CS_RNO[4]  (.A(\scalestate_0/N_1219 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO_1[4] ));
    NOR3A \scalestate_0/ACQ90_NUM_1_sqmuxa_0_a2_0  (.A(
        top_code_0_scaleload), .B(\top_code_0_scalechoice_0[4] ), .C(
        \top_code_0_scalechoice_0[1] ), .Y(\scalestate_0/N_62 ));
    XA1 \DUMP_OFF_1/off_on_timer_0/count_RNO[4]  (.A(
        \DUMP_OFF_1/off_on_timer_0/count_9_0 ), .B(
        \DUMP_OFF_1/count_4[4] ), .C(
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_n4 ));
    OR2B \top_code_0/n_acqnum_1_sqmuxa_0_o2  (.A(\xa_c[0] ), .B(
        \xa_c[1] ), .Y(\top_code_0/N_157 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m206  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[9] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_207 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[9]  (.A(
        \scalestate_0_strippluse[9] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[9] ));
    NOR2B \sd_acq_top_0/sd_sacq_state_0/cs_RNO[13]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_201 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[13] ));
    NOR2A \DDS_0/dds_state_0/w_clk_reg_RNIEMPL_0  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/w_clk_reg_net_1 ), .Y(
        \DDS_0/dds_state_0/para_1_sqmuxa_1 ));
    AO1 \state_1ms_0/timecount_RNO_2[15]  (.A(
        \state_1ms_0/M_DUMPTIME[15]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[15] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[15] ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg_RNI9SSG[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[0]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_0 ));
    OR3 \scalestate_0/timecount_ret_38_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[3] ), .B(
        \scalestate_0/OPENTIME_TEL_m[3] ), .C(
        \scalestate_0/timecount_20_iv_4[3] ), .Y(
        \scalestate_0/timecount_20_iv_8[3] ));
    DFN1E0 \DDS_0/dds_state_0/para[18]  (.D(\DDS_0/dds_state_0/N_163 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[18]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[4]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIABVJ2[13]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_1[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_0[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_12[0] ));
    MX2 \scalestate_0/dds_conf_RNO_0  (.A(\scalestate_0/un1_CS_20 ), 
        .B(scalestate_0_dds_conf), .S(\scalestate_0/N_1173 ), .Y(
        \scalestate_0/N_728 ));
    OR3 \scalestate_0/timecount_ret_54_RNIJ4I  (.A(
        \scalestate_0/timecount_20_0_iv_0_reto[19] ), .B(
        \scalestate_0/OPENTIME_TEL_m_reto[19] ), .C(
        \scalestate_0/timecount_20_0_iv_4_reto[19] ), .Y(
        \scalestate_0_timecount[19] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[13]_net_1 ));
    OR2 OR2_0 (.A(DUMP_0_dump_on), .B(DUMP_ON_0_dump_on), .Y(dumpon_c));
    DFN1 \timer_top_0/timer_0/timedata[9]  (.D(
        \timer_top_0/timer_0/timedata_4[9] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[9]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[5]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[5]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[5] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_52_i ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIGN2O3[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_7[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_18[0] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIMRJD[3]  (.A(
        \sd_acq_top_0/count_10[3] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[3]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_0[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_7[0] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIFAF91[2]  (.A(
        \ClockManagement_0/long_timer_0/count_c1 ), .B(
        \ClockManagement_0/long_timer_0/count[2]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c2 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_23  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[3] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[4] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[0] )
        );
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_1  (.A(
        \timer_top_0/dataout[6] ), .B(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_1_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_22[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[10]_net_1 ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_10[0] ));
    NOR2B \scalestate_0/s_acq180_RNO  (.A(\scalestate_0/N_742 ), .B(
        top_code_0_scale_rst), .Y(\scalestate_0/s_acq180_RNO_net_1 ));
    NOR2 \scalestate_0/M_NUM_1_sqmuxa_0_a2_0  (.A(
        \top_code_0_scalechoice_0[3] ), .B(
        \top_code_0_scalechoice_0[2] ), .Y(\scalestate_0/N_61 ));
    OR3 \DUMP_0/dump_coder_0/para6_RNI0E3J2[2]  (.A(
        \DUMP_0/dump_coder_0/i_reg16_3[0] ), .B(
        \DUMP_0/dump_coder_0/i_reg16_4[0] ), .C(
        \DUMP_0/dump_coder_0/i_reg16_NE_3[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_7[0] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[4]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c2 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n4 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[1] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[3]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c2 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n3 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[29]  (.D(
        \top_code_0_dds_configdata[12] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[29]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[5]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[5] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m39  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i22_mux ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m39 ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_13  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        , .B(\s_acq_change_0_s_stripnum[3] ), .C(
        \s_acq_change_0_s_stripnum[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_9 ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(\Signal_Noise_Acq_0/noise_acq_0/n_rdclk )
        );
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[3]  (.D(
        \top_code_0_bri_datain[13] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para3[3] ));
    NOR2B \top_code_0/relay_on_RNO[3]  (.A(\top_code_0/N_812 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[3]_net_1 ));
    NOR2A \timer_top_0/state_switch_0/state_over_n_RNO_0  (.A(
        \timer_top_0/state_switch_0/N_296 ), .B(
        noisestate_0_state_over_n), .Y(
        \timer_top_0/state_switch_0/N_278 ));
    NOR2B \PLUSE_0/qq_coder_0/i_RNO[0]  (.A(\PLUSE_0/up ), .B(
        bri_dump_sw_0_reset_out), .Y(\PLUSE_0/qq_coder_0/i_RNO_7[0] ));
    DFN1E1 \bridge_div_0/dataall[3]  (.D(\bridge_div_0/dataall_1[3] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/dataall[3]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/SXOR2_17_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_21_net ), 
        .B(\sd_acq_top_0/count[21] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[21] ));
    MX2 \scalestate_0/strippluse_RNO_2[8]  (.A(
        \scalestate_0/STRIPNUM180_NUM[8]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[8]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_428 ));
    DFN1 \timer_top_0/timer_0/timedata[13]  (.D(
        \timer_top_0/timer_0/timedata_4[13] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[13]_net_1 ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m46_5 ));
    IOPAD_TRI \GLA_pad/U0/U0  (.D(\GLA_pad/U0/NET1 ), .E(
        \GLA_pad/U0/NET2 ), .PAD(GLA));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[7]  (.A(
        \noisestate_0_timecount[7] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_205 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[5]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[5] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m124  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[3] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_125 ));
    NOR2B \top_code_0/plusedata_1_sqmuxa_0_a2_0_0  (.A(
        \top_code_0/N_340 ), .B(net_27), .Y(
        \top_code_0/plusedata_1_sqmuxa_0_a2_0_net_1 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[15]  (.A(\s_acq_change_0/N_85 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[15]_net_1 ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n5 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        );
    NOR3C \timer_top_0/timer_0/timedata_RNO[16]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_46 ), .Y(
        \timer_top_0/timer_0/timedata_4[16] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m239  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_240 ));
    NOR2A \GPMI_0/tri_state_0/xd_1  (.A(tri_ctrl_c), .B(zcs2_c), .Y(
        \GPMI_0.tri_state_0.xd_1 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_5_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/count_10[3] ), .C(\sd_acq_top_0/count_10[4] ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_5_net ));
    XOR2 \DUMP_0/dump_coder_0/para4_RNID82L[11]  (.A(
        \DUMP_0/dump_coder_0/para4[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_1_11[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m108  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[4] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_109 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[0]_net_1 ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n14 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        );
    IOTRI_OB_EB \s_acq180_pad/U0/U1  (.D(s_acq180_c), .E(VCC), .DOUT(
        \s_acq180_pad/U0/NET1 ), .EOUT(\s_acq180_pad/U0/NET2 ));
    OA1 \scalestate_0/timecount_ret_13_RNO  (.A(\scalestate_0/N_1267 ), 
        .B(\scalestate_0/N_1197 ), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/timecount_cnst_m_0[9] ));
    IOTRI_OB_EB \relay_on_pad[6]/U0/U1  (.D(\relay_on_c[6] ), .E(VCC), 
        .DOUT(\relay_on_pad[6]/U0/NET1 ), .EOUT(
        \relay_on_pad[6]/U0/NET2 ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_4  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[9]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] )
        );
    XOR2 \CAL_0/cal_div_0/count_RNI09VJ[4]  (.A(
        \CAL_0/cal_div_0/count[4]_net_1 ), .B(\CAL_0/cal_para_out[4] ), 
        .Y(\CAL_0/cal_div_0/clear_n4_4 ));
    NOR2B \scalestate_0/timecount_20_iv_4_RNO[5]  (.A(
        \scalestate_0/CUTTIMEI90[5]_net_1 ), .B(\scalestate_0/N_252 ), 
        .Y(\scalestate_0/CUTTIMEI90_m[5] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI3CQK[14]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[14]_net_1 ), .B(
        \sd_acq_top_0/count_0[14] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_14[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m176  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_177 ));
    NOR2 \PLUSE_0/qq_state_1/cs_RNO_1[3]  (.A(\PLUSE_0/i_2[2] ), .B(
        \PLUSE_0/qq_state_1/cs[3]_net_1 ), .Y(
        \PLUSE_0/qq_state_1/N_87 ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg_RNIKQP11[1]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[1]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_0 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[9]_net_1 ));
    DFN1 \scalestate_0/strippluse[6]  (.D(
        \scalestate_0/strippluse_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[6] ));
    DFN1E0 \DDS_0/dds_state_0/para[16]  (.D(\DDS_0/dds_state_0/N_18 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[16]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m263  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_260 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_263 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_264 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i10_mux ));
    AO1 \scalestate_0/necount_cmp_0/AO1_0  (.A(
        \scalestate_0/necount_cmp_0/AND2_0_Y ), .B(
        \scalestate_0/necount_cmp_0/NAND3A_1_Y ), .C(
        \scalestate_0/necount_cmp_0/NOR3_0_Y ), .Y(
        \scalestate_0/necount_cmp_0/AO1_0_Y ));
    DFN1E1 \plusestate_0/PLUSETIME[0]  (.D(\top_code_0_plusedata[0] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[0]_net_1 ));
    NOR2B \DSTimer_0/dump_sustain_timer_0/data_RNO[1]  (.A(
        \DSTimer_0/dump_sustain_timer_0/N_25 ), .B(
        top_code_0_dump_sustain), .Y(
        \DSTimer_0/dump_sustain_timer_0/data_RNO[1]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[15]  (.A(
        \state_1ms_0/PLUSECYCLE[15]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[15] ));
    NOR2B \scalestate_0/timecount_RNO_1[20]  (.A(
        \scalestate_0/OPENTIME_TEL[20]_net_1 ), .B(
        \scalestate_0/N_258 ), .Y(\scalestate_0/OPENTIME_TEL_m[20] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m32  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_31 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_32 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_33 ));
    XOR2 \scalestate_0/M_pulse_RNO_5  (.A(
        \scalestate_0/M_NUM[10]_net_1 ), .B(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/M_pulse8_10 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_11_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_154_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_58_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_11_inst ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/OAND2_24_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net ), 
        .C(\sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_19_net ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[3] ));
    DFN1 \nsctrl_choice_0/dumponoff_rst  (.D(
        \nsctrl_choice_0/dumponoff_rst_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(nsctrl_choice_0_dumponoff_rst));
    AND2 \ClockManagement_0/clk_div500_0/un1_count_1_I_1  (.A(
        \ClockManagement_0/clk_div500_0/count[0]_net_1 ), .B(
        \ClockManagement_0/clk_5M_en ), .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_TMP[0] ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[2]_net_1 ));
    DFN1 \scalestate_0/reset_out  (.D(
        \scalestate_0/reset_out_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        net_45));
    NOR2B \DDS_0/dds_coder_0/i_RNO_1[3]  (.A(\DDS_0/count[6] ), .B(
        \DDS_0/count[5] ), .Y(\DDS_0/dds_coder_0/m8_1 ));
    OAI1 \plusestate_0/timecount_1_RNO_1[7]  (.A(
        \plusestate_0/CS[4]_net_1 ), .B(\plusestate_0/CS[8]_net_1 ), 
        .C(top_code_0_pluse_rst_0), .Y(\plusestate_0/N_253 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m45_2 ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_1_Y ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_19  (.A(
        \timer_top_0/dataout[15] ), .B(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_19_Y ));
    DFN1E1 \scalestate_0/timecount_ret_46  (.D(
        \scalestate_0/OPENTIME_TEL_m[16] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/OPENTIME_TEL_m_reto[16] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[4]  (.A(
        \scalestate_0_timecount[4] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_223 ));
    NOR2B \sd_acq_top_0/sd_sacq_state_0/cs_RNO[7]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_203 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[7] ));
    MX2 \top_code_0/relay_close_RNO_0[9]  (.A(\relay_close_c[9] ), .B(
        \GPMI_0_dataout[9] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_828 ));
    DFN1E1 \scalestate_0/CUTTIME90[7]  (.D(\top_code_0_scaledatain[7] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[7]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m286  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_283 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_286 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_287 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNITVDS[12]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[12]_net_1 ), .B(
        \sd_acq_top_0/count_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_12[0] ));
    XA1 \DDS_0/dds_timer_0/count_RNO[4]  (.A(
        \DDS_0/dds_timer_0/count_c3 ), .B(\DDS_0/count[4] ), .C(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DDS_0/dds_timer_0/count_n4 ));
    OA1B \syn_md_module_1/syn_md_0/count_RNO[1]  (.A(
        \syn_md_module_1/syn_md_0/N_23_1 ), .B(
        \syn_md_module_1/syn_md_0/count_RNO_0[1]_net_1 ), .C(
        \syn_md_module_1/syn_md_0/N_50 ), .Y(
        \syn_md_module_1/syn_md_0/count_RNO[1]_net_1 ));
    IOBI_IB_OB_EB \xd_pad[11]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[11] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[11]/U0/NET3 ), .DOUT(
        \xd_pad[11]/U0/NET1 ), .EOUT(\xd_pad[11]/U0/NET2 ), .Y(
        \xd_in[11] ));
    OR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_4  (
        .A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[4]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_5 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_6  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_146_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_100_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_6_Y ));
    DFN1 \top_code_0/scan_rst_0_0  (.D(
        \top_code_0/scan_rst_RNIMNCI3_net_1 ), .CLK(GLA_net_1), .Q(
        net_33_0));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIPRDS[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[10]_net_1 ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_10[0] ));
    OR3 \scalestate_0/timecount_ret_82_RNO  (.A(
        \scalestate_0/PLUSETIME90_m[4] ), .B(
        \scalestate_0/DUMPTIME_m[4] ), .C(
        \scalestate_0/S_DUMPTIME_m[4] ), .Y(
        \scalestate_0/timecount_20_iv_6[4] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_103  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_59_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_120_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_103_Y ));
    DFN1 \DUMP_0/dump_timer_0/count[9]  (.D(
        \DUMP_0/dump_timer_0/count_n9 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count[9] ));
    MX2 \scalestate_0/strippluse_RNO_0[3]  (.A(
        \scalestate_0/strippluse_6[3] ), .B(
        \scalestate_0_strippluse[3] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_562 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[28]  (.A(
        \top_code_0_dds_configdata[11] ), .B(\DDS_0/dds_state_0/N_569 )
        , .C(\DDS_0/dds_state_0/N_478 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[28] ));
    DFN1 \ClockManagement_0/clk_div500_0/count[7]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[7] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[7]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_6[14]  (.A(
        \state_1ms_0/PLUSETIME[14]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[14] ));
    NOR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en_net_1 ), .B(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_6 ));
    OAI1 \scalestate_0/CS_RNI96JS[5]  (.A(scalestate_0_ne_le), .B(
        \scalestate_0/CS[5]_net_1 ), .C(top_code_0_scale_rst_3), .Y(
        \scalestate_0/timecount_8_sqmuxa_i_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_54_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_60  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_60_Y ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[2] ), .CLK(
        GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[12]  (.A(
        \noisestate_0/acqtime[12]_net_1 ), .B(
        \noisestate_0/dectime[12]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_69 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i8_mux ));
    AO1 \state_1ms_0/timecount_RNO_4[8]  (.A(
        \state_1ms_0/S_DUMPTIME[8]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[8] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[8] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[6]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[5]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c4 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n6 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[8]  (.A(
        \timer_top_0/state_switch_0/N_245 ), .B(
        \timer_top_0/state_switch_0/N_246 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[8] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[8]_net_1 ));
    DFN1 \PLUSE_0/qq_state_0/cs[3]  (.D(
        \PLUSE_0/qq_state_0/cs_RNO_1[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/qq_state_0/cs[3]_net_1 ));
    NOR2B \DDS_0/dds_state_0/w_clk_RNO  (.A(
        \DDS_0/dds_state_0/w_clk_reg_net_1 ), .B(
        \DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/w_clk_RNO_net_1 ));
    XOR2 \ClockManagement_0/clk_div500_0/un1_count_1_I_35  (.A(
        \ClockManagement_0/clk_div500_0/count[2]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_1[0] ), 
        .Y(\ClockManagement_0/clk_div500_0/I_35 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[8]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n8 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ));
    DFN1 \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1  (.D(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(\GPMI_0/xwe_xzcs2_syn_0/xwe_reg1_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[20]  (.A(
        \top_code_0_dds_configdata[3] ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_466 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[20] ));
    DFN1E1 \top_code_0/scandata[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[1] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_45  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_45_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_49  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_1_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_1_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_49_Y ));
    OR3A \top_code_0/n_rd_en_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/N_207 ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_17  (.A(\PLUSE_0/count_8[4] ), 
        .B(\PLUSE_0/half_para[4] ), .Y(\PLUSE_0/bri_coder_0/N_5 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[8]  (.D(
        \top_code_0_dds_configdata[7] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[8]_net_1 ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[4]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_31 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[4] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNILCUE[1]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[1]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_1[0] ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[2]_net_1 ));
    DFN1E1 \noisestate_0/dectime[0]  (.D(\top_code_0_noisedata[0] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[0]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m44_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[15] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[2]  (.D(
        \top_code_0_pd_pluse_data[2] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[2]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m188  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_185 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_188 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_189 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[0]  (.A(
        \scalestate_0_timecount[0] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_243 ));
    IOTRI_OB_EB \relay_on_pad[0]/U0/U1  (.D(\relay_on_c[0] ), .E(VCC), 
        .DOUT(\relay_on_pad[0]/U0/NET1 ), .EOUT(
        \relay_on_pad[0]/U0/NET2 ));
    XA1 \DUMP_0/off_on_timer_0/count_RNO[4]  (.A(
        \DUMP_0/off_on_timer_0/count_9_0 ), .B(\DUMP_0/count_2[4] ), 
        .C(\DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_0/count_n4 ));
    NOR3A \scalestate_0/necount_cmp_1/NOR3A_1  (.A(
        \scalestate_0/necount_cmp_1/OR2A_2_Y ), .B(
        \scalestate_0/necount_cmp_1/AO1C_1_Y ), .C(
        \scalestate_0/NE_NUM[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/NOR3A_1_Y ));
    OR3A \top_code_0/RAM_Rd_rst_3_i_o2_0  (.A(\xa_c[4] ), .B(
        \top_code_0/N_139 ), .C(\xa_c[7] ), .Y(\top_code_0/N_155 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[11]  (.D(
        \top_code_0_state_1ms_data[11] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[11]_net_1 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[4]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_4[4] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[4]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_84  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_45_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_56_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_84_Y ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[8]  (.A(
        \DUMP_0/dump_timer_0/count_c7 ), .B(\DUMP_0/count[8] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n8 ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_6_inst  (.A(
        \scalestate_0/necount_inc_0/Rcout_8_net ), .B(
        \scalestate_0/necount[8]_net_1 ), .Y(
        \scalestate_0/necount1[8] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[10] ));
    NOR2B \state_1ms_0/timecount_RNO_6[12]  (.A(
        \state_1ms_0/PLUSETIME[12]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[12] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[6]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[6] ));
    DFN1E1 \top_code_0/s_addchoice_2[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_2[4] ));
    DFN1E1 \scalestate_0/OPENTIME[6]  (.D(\top_code_0_scaledatain[6] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[6]_net_1 ));
    NOR3A \DUMP_0/dump_state_0/un1_ns_0_a2  (.A(\DUMP_0/i[8] ), .B(
        \DUMP_0/i[6] ), .C(\DUMP_0/i[4] ), .Y(
        \DUMP_0/dump_state_0/N_201 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[8] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[1]  (.D(
        \top_code_0_halfdata_0[1] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[1] ));
    NOR2B \DUMP_0/dump_coder_0/para18  (.A(\top_code_0_dump_cho_0[0] ), 
        .B(\top_code_0_dump_cho_0[1] ), .Y(
        \DUMP_0/dump_coder_0/para18_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m259  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_258 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_259 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_260 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[9] ));
    AND2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/QAND2_25_inst  (
        .A(\sd_acq_top_0/count[18] ), .B(\sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_31_net ));
    OR3 \top_code_0/pn_change_RNO_0  (.A(\top_code_0/N_144 ), .B(
        \top_code_0/N_148 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/N_219 ));
    AO1A \scanstate_0/dds_conf_RNO_0  (.A(\scanstate_0/CS[2]_net_1 ), 
        .B(scanstate_0_dds_conf), .C(\scanstate_0/CS[1]_net_1 ), .Y(
        \scanstate_0/N_130 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[13]_net_1 ));
    AND3 \scalestate_0/necount_cmp_0/AND3_0  (.A(
        \scalestate_0/necount_cmp_0/AND3_1_Y ), .B(
        \scalestate_0/necount_cmp_0/XNOR2_6_Y ), .C(
        \scalestate_0/necount_cmp_0/XNOR2_4_Y ), .Y(
        \scalestate_0/necount_cmp_0/AND3_0_Y ));
    DFN1E1 \scalestate_0/timecount_ret_66  (.D(
        \scalestate_0/timecount_20_iv_7[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[14] ));
    NOR3A \dds_change_0/dds_conf_RNO_4  (.A(scanstate_0_dds_conf), .B(
        \top_code_0_change_0[0] ), .C(\top_code_0_change_0[1] ), .Y(
        \dds_change_0/dds_confin1_m ));
    IOTRI_OB_EB \relay_close_pad[7]/U0/U1  (.D(\relay_close_c[7] ), .E(
        VCC), .DOUT(\relay_close_pad[7]/U0/NET1 ), .EOUT(
        \relay_close_pad[7]/U0/NET2 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m16  
        (.A(\s_acq_change_0_s_stripnum[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[5]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i10_mux )
        );
    OA1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[3]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/en1 ), .B(\sd_acq_top_0/i_1[5] ), 
        .C(\sd_acq_top_0/sd_sacq_state_0/cs[2]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_237 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[2]  (.D(
        \top_code_0_n_divnum_0[2] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[2]_net_1 ));
    DFN1 \scalestate_0/pluse_start  (.D(
        \scalestate_0/pluse_start_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_pluse_start));
    NOR2A \s_acq_change_0/s_acqnum_RNO_1[12]  (.A(
        \top_code_0_s_acqnum_2[12] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[12] ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI4S898[1]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_11[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_10[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_12[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_i[0] ));
    XA1C \DUMP_0/dump_coder_0/i_RNO_5[3]  (.A(\DUMP_0/count_1[4] ), .B(
        \DUMP_0/dump_coder_0/para1[4]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_5[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_3[3] ));
    NOR2 \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[3]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/en1 ), .B(\sd_acq_top_0/i_2[4] ), 
        .Y(\sd_acq_top_0/sd_sacq_state_0/N_236 ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_7  (.A(
        \scalestate_0/NE_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_7_Y ));
    DFN1 \PLUSE_0/qq_timer_1/count[4]  (.D(
        \PLUSE_0/qq_timer_1/count_n4 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_7[4] ));
    IOBI_IB_OB_EB \xd_pad[8]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[8] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[8]/U0/NET3 ), .DOUT(\xd_pad[8]/U0/NET1 ), .EOUT(
        \xd_pad[8]/U0/NET2 ), .Y(\xd_in[8] ));
    DFN1 \bri_dump_sw_0/reset_out_0_0  (.D(
        \bri_dump_sw_0/reset_out_0_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_reset_out_0));
    DFN1E1 \state_1ms_0/CUTTIME[3]  (.D(\top_code_0_state_1ms_data[3] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[3]_net_1 ));
    NOR3 \top_code_0/sigrst_RNO_1  (.A(\top_code_0/N_151 ), .B(
        \top_code_0/N_158 ), .C(\top_code_0/N_159 ), .Y(
        \top_code_0/N_312 ));
    AND3 \scalestate_0/necount_inc_0/AND2_9_inst  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .C(
        \scalestate_0/necount[8]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/inc_10_net ));
    NOR3 \top_code_0/un1_xa_2_0_a2_1  (.A(\xa_c[18] ), .B(
        \top_code_0/un1_xa_30_0_o2_0_net_1 ), .C(\xa_c[6] ), .Y(
        \top_code_0/N_336 ));
    DFN1E1 \top_code_0/state_1ms_data[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[1] ));
    DFN1E1 \top_code_0/dumpdata[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[8] ));
    DFN1E1 \scalestate_0/OPENTIME[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[15]_net_1 ));
    XOR2 \PLUSE_0/qq_coder_0/i_reg10_3[0]  (.A(\PLUSE_0/qq_para3[3] ), 
        .B(\PLUSE_0/count_9[3] ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_3[0]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m234  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_227 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_234 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[8] ));
    DFN1 \nsctrl_choice_0/soft_d  (.D(
        \nsctrl_choice_0/soft_d_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_soft_d));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_48  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_50_i ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[6] )
        );
    NAND3A \scalestate_0/necount_cmp_1/NAND3A_2  (.A(
        \scalestate_0/NE_NUM[4]_net_1 ), .B(
        \scalestate_0/necount[4]_net_1 ), .C(
        \scalestate_0/necount_cmp_1/OR2A_0_Y ), .Y(
        \scalestate_0/necount_cmp_1/NAND3A_2_Y ));
    IOBI_IB_OB_EB \xd_pad[12]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[12] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[12]/U0/NET3 ), .DOUT(
        \xd_pad[12]/U0/NET1 ), .EOUT(\xd_pad[12]/U0/NET2 ), .Y(
        \xd_in[12] ));
    MX2 \top_code_0/relay_close_RNO_0[4]  (.A(\relay_close_c[4] ), .B(
        \GPMI_0_dataout[4] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_823 ));
    DFN1 \timer_top_0/state_switch_0/clk_en_noise  (.D(
        \timer_top_0/state_switch_0/clk_en_noise_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(timer_top_0_clk_en_noise));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[13]  (.A(
        \timer_top_0/state_switch_0/N_190 ), .B(
        \timer_top_0/state_switch_0/N_191 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[13] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[13]_net_1 ));
    OR3 \scalestate_0/timecount_ret_66_RNIS7I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[14] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[14] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[14] ), .Y(
        \scalestate_0_timecount[14] ));
    NOR3B \PLUSE_0/bri_timer_0/clken  (.A(pulse_start_c), .B(clk_4f_en)
        , .C(\PLUSE_0/bri_coder_0_half ), .Y(
        \PLUSE_0/bri_timer_0/clken_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIS7811[13]  (.A(
        \sd_acq_top_0/count_0[13] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[13]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_11[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_1[0] ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[13]  (.A(
        \ClockManagement_0/long_timer_0/count_c12 ), .B(
        \ClockManagement_0/long_timer_0/count[13]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n13 ));
    AO1 \timer_top_0/state_switch_0/dataout_RNO[17]  (.A(
        \state_1ms_0_timecount[17] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .C(
        \timer_top_0/state_switch_0/N_268 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[17]_net_1 ));
    DFN1 \top_code_0/scale_rst  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[1]  (.A(
        \plusestate_0_timecount[1] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_239 ));
    NOR2A \scalestate_0/timecount_ret_85_RNO_1  (.A(
        \scalestate_0/DUMPTIME[11]_net_1 ), .B(\scalestate_0/N_1093 ), 
        .Y(\scalestate_0/DUMPTIME_m[11] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[26]  (.A(
        \top_code_0_dds_configdata[9] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_470 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[26] ));
    NOR2A \state_1ms_0/timecount_RNO_5[6]  (.A(
        \state_1ms_0/CS[5]_net_1 ), .B(
        \state_1ms_0/PLUSETIME[6]_net_1 ), .Y(
        \state_1ms_0/PLUSETIME_i_m[6] ));
    MX2 \PLUSE_0/bri_timer_0/count[6]/U0  (.A(\PLUSE_0/count_2[6] ), 
        .B(\PLUSE_0/bri_timer_0/count_n6 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[6]/Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m217  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_216 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_217 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_218 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m70  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m70_4 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[2] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_4  (.A(\ADC_c[6] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ));
    AND2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_8  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[1] )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m146  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_145 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_146 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_147 ));
    OR3A \top_code_0/dds_load_RNO_0  (.A(\xa_c[1] ), .B(
        \top_code_0/N_142 ), .C(\top_code_0/N_155 ), .Y(
        \top_code_0/N_200 ));
    MX2 \noisestate_0/timecount_1_RNO_0[14]  (.A(
        \noisestate_0/acqtime[14]_net_1 ), .B(
        \noisestate_0/dectime[14]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_71 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[0]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1[0] ), 
        .CLK(GLA_net_1), .E(top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[0]_net_1 ));
    XA1C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_10[4]  (.A(
        \pd_pluse_top_0/count_0[8] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[8]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_13[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_2[4] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[2]  (.A(
        \scalestate_0/s_acqnum_7[2] ), .B(\scalestate_0_s_acqnum[2] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_549 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[3]  (.A(
        \top_code_0_dumpdata_0[3] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[3] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m61  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[16] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_62 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i10_mux ));
    MX2 \scalestate_0/CS_RNO_0[4]  (.A(\scalestate_0/CS[4]_net_1 ), .B(
        \scalestate_0/CS[19]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1219 ));
    OR2A \noisestate_0/CS_RNI1M6C[6]  (.A(top_code_0_noise_rst), .B(
        \noisestate_0/N_250 ), .Y(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I10_un1_CO1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N168 ), 
        .B(\s_acq_change_0_s_stripnum[10] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I10_un1_CO1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIQ009[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[0]_net_1 ), .B(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_0[0] ));
    MX2B \PLUSE_0/bri_state_0/cs_RNO[14]  (.A(
        \PLUSE_0/bri_state_0/cs[14]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[13] ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_RNO[14]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m45_4 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_9[3]  (.A(
        \DUMP_0/dump_coder_0/para1[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_10[0] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[3]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c2 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n3 ));
    AO1C \scanstate_0/CS_RNO_0[2]  (.A(\scanstate_0/CS[1]_net_1 ), .B(
        timer_top_0_clk_en_scan), .C(net_33_0), .Y(
        \scanstate_0/CS_srsts_i_0[2] ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[2]  (.A(\s_acq_change_0/N_72 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[2]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m45  
        (.A(\s_acq_change_0_s_stripnum[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[9]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i16_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_46_i ));
    MX2 \nsctrl_choice_0/dumpoff_ctr_RNO_0  (.A(
        scanstate_0_dumpoff_ctr), .B(noisestate_0_dumpoff_ctr), .S(
        top_code_0_n_s_ctrl_1), .Y(\nsctrl_choice_0/dumpoff_ctr_5 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIMRID1[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_3[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_10[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_7[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_11[0] ));
    DFN1E1 \top_code_0/scaledatain[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[15] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[11]  (.A(
        \scanstate_0_timecount[11] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_196 ));
    NOR2B \scanstate_0/dds_conf_RNO  (.A(\scanstate_0/N_130 ), .B(
        net_33), .Y(\scanstate_0/dds_conf_RNO_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[1]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[1] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[1] ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[3]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[3] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_10[3] ));
    AND2A \scalestate_0/necount_cmp_1/AND2A_0  (.A(
        \scalestate_0/necount[10]_net_1 ), .B(
        \scalestate_0/NE_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/AND2A_0_Y ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[0]  (.D(
        \top_code_0_pd_pluse_data[0] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[0]_net_1 ));
    AX1C \bridge_div_0/count_5_I_12  (.A(
        \bridge_div_0/count_RNIHPOM7[3]_net_1 ), .B(
        \bridge_div_0/DWACT_FINC_E[0] ), .C(
        \bridge_div_0/count_RNIIQOM7[4]_net_1 ), .Y(
        \bridge_div_0/count_5[4] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_58_i ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m17  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_16_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_17_0 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_18_0 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIKE6P1[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_11[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_13[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_13[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m306  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[12] ), .C(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_307 ));
    NOR2A \scalestate_0/timecount_ret_33_RNO_0  (.A(
        \scalestate_0/timecount_cnst[1] ), .B(\scalestate_0/N_258_0 ), 
        .Y(\scalestate_0/timecount_m1_e_2_0 ));
    MX2 \noisestate_0/sw_acq2_RNO_0  (.A(noisestate_0_sw_acq2), .B(
        \noisestate_0/N_233 ), .S(\noisestate_0/N_248 ), .Y(
        \noisestate_0/N_108 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[11]  (.A(
        \ClockManagement_0/long_timer_0/count_c10 ), .B(
        \ClockManagement_0/long_timer_0/count[11]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n11 ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_7  (.A(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .B(
        \timer_top_0/dataout[7] ), .C(
        \timer_top_0/timer_0/timedata[6]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_7_Y ));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[5]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_187 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_176 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_2[5] ));
    DFN1E1 \top_code_0/bri_datain[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[3] ));
    DFN1 \noisestate_0/CS_i_0[0]  (.D(
        \noisestate_0/CS_i_0_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \noisestate_0/CS_li[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m107  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_106 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_107 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_108 ));
    OR3 \scalestate_0/timecount_ret_77_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[6] ), .B(
        \scalestate_0/OPENTIME_TEL_m[6] ), .C(
        \scalestate_0/timecount_20_iv_4[6] ), .Y(
        \scalestate_0/timecount_20_iv_8[6] ));
    NOR2A \scalestate_0/necount_LE_NE_RNIQ3SG  (.A(
        \scalestate_0/CS[11]_net_1 ), .B(scalestate_0_ne_le), .Y(
        \scalestate_0/N_1267 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[2]  (.A(
        \scalestate_0_strippluse[2] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[2] ));
    IOPAD_TRI \rt_sw_pad/U0/U0  (.D(\rt_sw_pad/U0/NET1 ), .E(
        \rt_sw_pad/U0/NET2 ), .PAD(rt_sw));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[9]  (.A(
        \noisestate_0_timecount[9] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_200 ));
    DFN1 \syn_md_module_1/syn_md_0/count[1]  (.D(
        \syn_md_module_1/syn_md_0/count_RNO[1]_net_1 ), .CLK(GLA_net_1)
        , .Q(\syn_md_module_1/syn_md_0/count[1]_net_1 ));
    OR3 \DUMP_0/dump_coder_0/para4_RNICE047[10]  (.A(
        \DUMP_0/dump_coder_0/un1_count_1_NE_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_NE_6[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_1_NE_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_108  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_132_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_82_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_108_Y ));
    NOR2A \DUMP_0/dump_state_0/cs_RNO_1[2]  (.A(\DUMP_0/i_0[2] ), .B(
        \DUMP_0/dump_state_0/cs[1]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_183 ));
    OR2A \top_code_0/noise_rst_0_0_RNIDOO43  (.A(net_27), .B(
        \top_code_0/N_805 ), .Y(
        \top_code_0/noise_rst_0_0_RNIDOO43_net_1 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNISCF21[10]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_4 ), .B(
        \s_acq_change_0_s_stripnum[10] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_10 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_12  (.A(
        \timer_top_0/dataout[13] ), .B(
        \timer_top_0/timer_0/timedata[13]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_12_Y ));
    DFN1 \s_acq_change_0/s_stripnum[5]  (.D(
        \s_acq_change_0/s_stripnum_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[5] ));
    DFN1 \scan_scale_sw_0/s_start  (.D(
        \scan_scale_sw_0/s_start_RNO_net_1 ), .CLK(ddsclkout_c), .Q(
        scan_scale_sw_0_s_start));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_38  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_52_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[1] )
        );
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m175  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_176 ));
    OA1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_11  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_11 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_11 ));
    OR3 \scalestate_0/timecount_ret_22_RNIO7I  (.A(
        \scalestate_0/timecount_20_iv_3_reto[10] ), .B(
        \scalestate_0/timecount_20_iv_2_reto[10] ), .C(
        \scalestate_0/timecount_20_iv_6_reto[10] ), .Y(
        \scalestate_0/timecount_20_iv_9_reto[10] ));
    NOR2B \top_code_0/relay_on_RNO[4]  (.A(\top_code_0/N_813 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[4]_net_1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[11]  (.A(
        \s_acq_change_0/s_stripnum_5[11] ), .B(
        \s_acq_change_0_s_stripnum[11] ), .S(\top_code_0_change[1] ), 
        .Y(\s_acq_change_0/N_67 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[12]  (.D(
        \top_code_0_pd_pluse_data[12] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[12]_net_1 ));
    NOR2B \top_code_0/noisedata_1_sqmuxa_0_a2_0  (.A(\xa_c[3] ), .B(
        \top_code_0/N_329 ), .Y(\top_code_0/N_333 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m21  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_22 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/ADD_20x20_slow_I19_Y_3 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[19] ));
    XA1 \DSTimer_0/dump_sustain_timer_0/count_RNO[3]  (.A(
        \DSTimer_0/dump_sustain_timer_0/count_7_0 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[3]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p ), .Y(
        \DSTimer_0/dump_sustain_timer_0/count_n3 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[4]  (.A(\DDS_0/dds_state_0/N_318 )
        , .B(\DDS_0/dds_state_0/N_317 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[4] ), .Y(
        \DDS_0/dds_state_0/N_54 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[17]  (.A(
        \DDS_0/dds_state_0/N_500 ), .B(\DDS_0/dds_state_0/N_499 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[17] ), .Y(
        \DDS_0/dds_state_0/N_161 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[13]  (.A(
        \DDS_0/dds_state_0/N_337 ), .B(\DDS_0/dds_state_0/N_336 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[13] ), .Y(
        \DDS_0/dds_state_0/N_118 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[7]_net_1 ));
    DFN1E1 \top_code_0/pd_pluse_data[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[13] ));
    DFN1E0 \DDS_0/dds_state_0/para[25]  (.D(\DDS_0/dds_state_0/N_25 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[25]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_41_RNO_4  (.A(
        \scalestate_0/CUTTIMEI90[2]_net_1 ), .B(\scalestate_0/N_252 ), 
        .Y(\scalestate_0/CUTTIMEI90_m[2] ));
    NOR2B \DUMP_0/dump_state_0/cs_RNIRPGC[5]  (.A(
        \DUMP_0/dump_state_0_on_start ), .B(
        \DUMP_0/dump_state_0/N_206 ), .Y(
        \DUMP_0/dump_state_0/un1_ns_0_a3_0 ));
    OA1 \pd_pluse_top_0/pd_pluse_state_0/en_RNO  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/en2 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/en1_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/en_RNO_net_1 ));
    DFN1E1 \top_code_0/pd_pluse_choice[0]  (.D(\GPMI_0_dataout[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_choice_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_choice[0] ));
    MX2A \scalestate_0/fst_lst_pulse_RNO_0  (.A(
        \scalestate_0/fst_lst_pulse8_NE ), .B(
        \scalestate_0/fst_lst_pulse_net_1 ), .S(\scalestate_0/N_1181 ), 
        .Y(\scalestate_0/N_741 ));
    AO1C \scanstate_0/CS_RNO_0[5]  (.A(\scanstate_0/CS[4]_net_1 ), .B(
        timer_top_0_clk_en_scan), .C(net_33), .Y(
        \scanstate_0/CS_srsts_i_0[5] ));
    OAI1 \scalestate_0/dump_sustain_ctrl_RNO_1  (.A(
        \scalestate_0/CS_0[11]_net_1 ), .B(\scalestate_0/CS[13]_net_1 )
        , .C(timer_top_0_clk_en_scale_0), .Y(\scalestate_0/N_1183 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[11]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[11]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_327 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_10_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_10_net ));
    MX2 \scanstate_0/timecount_1_RNO_0[9]  (.A(
        \scanstate_0/dectime[9]_net_1 ), .B(
        \scanstate_0/acqtime[9]_net_1 ), .S(\scanstate_0/CS[4]_net_1 ), 
        .Y(\scanstate_0/N_67 ));
    OR3B \scalestate_0/timecount_ret_33_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS_i[0]_net_1 ), .C(
        \scalestate_0/un1_CS_20 ), .Y(\scalestate_0/timecount_cnst[1] )
        );
    XA1 \DUMP_0/off_on_timer_0/count_RNO[1]  (.A(\DUMP_0/count_2[1] ), 
        .B(\DUMP_0/count_2[0] ), .C(
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_0/count_n1 ));
    AO1A \scalestate_0/timecount_ret_70_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[15]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[15] ), .Y(
        \scalestate_0/timecount_20_iv_1[15] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_13  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_13_Y ));
    DFN1E0 \DDS_0/dds_state_0/para[21]  (.D(\DDS_0/dds_state_0/N_167 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[21]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m233  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_230 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_233 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_234 ));
    DFN1 \ClockManagement_0/clk_10k_0/clk_5M_reg2  (.D(
        \ClockManagement_0/clk_10k_0/clk_5M_reg2_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(\ClockManagement_0/clk_10k_0/clk_5M_reg2_net_1 )
        );
    OR3 \top_code_0/n_load_RNO_0  (.A(\top_code_0/N_154 ), .B(
        \top_code_0/N_152 ), .C(\top_code_0/N_147 ), .Y(
        \top_code_0/N_201 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNISJ0I1[12]  (.A(
        \sd_acq_top_0/count_0[12] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[12]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_7[0] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[2]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[2] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[20]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[20]_net_1 ));
    XNOR2 \PLUSE_0/bri_coder_0/half_0_I_2  (.A(\PLUSE_0/half_para[6] ), 
        .B(\PLUSE_0/count_2[6] ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[1] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIS5KE3[7]  (.A(
        \ClockManagement_0/long_timer_0/count_c6 ), .B(
        \ClockManagement_0/long_timer_0/count[7]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c7 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[9]  (.A(
        \state_1ms_0_timecount[9] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_202 ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIS0T91[15]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[14]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_0 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_7 ));
    DFN1E1 \scalestate_0/PLUSETIME90[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[0]_net_1 ));
    DFN1E1 \scalestate_0/ACQTIME[0]  (.D(\top_code_0_scaledatain_0[0] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[0]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_8[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[9]_net_1 ), .B(
        \pd_pluse_top_0/count_0[9] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_9[0] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_7  (.A(
        \timer_top_0/dataout[17] ), .B(
        \timer_top_0/timer_0/timedata[17]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_7_Y ));
    DFN1E1 \scalestate_0/DUMPTIME[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[11]_net_1 ));
    MX2 \top_code_0/relay_on_RNO_0[2]  (.A(\relay_on_c[2] ), .B(
        \GPMI_0_dataout[2] ), .S(\top_code_0/relay_on_1_sqmuxa ), .Y(
        \top_code_0/N_811 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI8C521[14]  (.A(
        \sd_acq_top_0/count_0[14] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[14]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_8[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_0[0] ));
    DFN1 \state_1ms_0/timecount[5]  (.D(
        \state_1ms_0/timecount_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[5] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_71  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_71_Y ));
    DFN1C0 \PLUSE_0/bri_state_0/up/U1  (.D(\PLUSE_0/bri_state_0/up/Y ), 
        .CLK(ddsclkout_c), .CLR(\PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/up ));
    NOR2A \scalestate_0/timecount_ret_59_RNO_4  (.A(
        \scalestate_0/CUTTIME90[0]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[0] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI6H6B[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_5[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m254  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[15] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_255 ));
    NOR2B \DUMP_OFF_0/off_on_timer_0/count_RNIPI3G[2]  (.A(
        \DUMP_OFF_0/off_on_timer_0/count_c1 ), .B(
        \DUMP_OFF_0/count_3[2] ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_c2 ));
    NOR2A \bridge_div_0/count_RNIQJF17[3]  (.A(
        \bridge_div_0/clear1_n17_NE[0] ), .B(
        \bridge_div_0/un1_count_i[0] ), .Y(\bridge_div_0/clear1_n18 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m300  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_299 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_300 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_301 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_1_net_1 )
        );
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[1]  (.D(
        \top_code_0_n_acqnum_2[1] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[1]_net_1 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[0]  (.D(\top_code_0_scaledatain[0] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[0]_net_1 ));
    IOPAD_IN \xa_pad[0]/U0/U0  (.PAD(xa[0]), .Y(\xa_pad[0]/U0/NET1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m215  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[9] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_216 ));
    DFN1E1 \top_code_0/plusedata[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[0] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[2]  (.A(\scalestate_0/N_450 ), 
        .B(\scalestate_0/ACQECHO_NUM[2]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[2] ));
    DFN1 \DSTimer_0/dump_sustain_timer_0/count[2]  (.D(
        \DSTimer_0/dump_sustain_timer_0/count_n2 ), .CLK(clock_10khz), 
        .Q(\DSTimer_0/dump_sustain_timer_0/count[2]_net_1 ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_9  (.A(\ADC_c[1] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_9 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[6]  (.D(\top_code_0_scaledatain[6] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[6]_net_1 ));
    OR3 \DUMP_0/dump_coder_0/para3_RNI4DB52[10]  (.A(
        \DUMP_0/dump_coder_0/un1_count_2_10[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_2_0_0[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_8[0] ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[3]  (.A(
        \s_acq_change_0/s_stripnum_5[3] ), .B(
        \s_acq_change_0_s_stripnum[3] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_59 ));
    XA1A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_9[10]  (.A(
        \sd_acq_top_0/count_10[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[0]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_11[10] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[5]  (.A(
        \scalestate_0_timecount[5] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_218 ));
    DFN1E1 \scalestate_0/PLUSETIME90[2]  (.D(
        \top_code_0_scaledatain[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[2]_net_1 ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_6  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/M_NUM[9]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_6_Y ));
    OR2 \top_code_0/bridge_load_3_i_o3  (.A(\top_code_0/N_174 ), .B(
        \top_code_0/N_157 ), .Y(\top_code_0/N_216 ));
    NOR3 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m4_e  (.A(
        \top_code_0_s_addchoice[2] ), .B(\top_code_0_s_addchoice[3] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_311 ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_313 ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_20  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[0] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[2] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[3] )
        );
    NOR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[5]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_216 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_217 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[5] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[11]  (.A(\scalestate_0/N_459 ), 
        .B(\scalestate_0/ACQECHO_NUM[11]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[11] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[19]  (.D(
        \top_code_0_dds_configdata[2] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[19]_net_1 ));
    OR2B \scalestate_0/CS_RNI8O8M[13]  (.A(\scalestate_0/CS[13]_net_1 )
        , .B(\scalestate_0/N_1196 ), .Y(\scalestate_0/N_1179 ));
    OR3 \syn_md_module_1/syn_md_0/count_RNII9OC[2]  (.A(
        \syn_md_module_1/syn_md_0/count[0]_net_1 ), .B(
        \syn_md_module_1/syn_md_0/count[1]_net_1 ), .C(
        \syn_md_module_1/syn_md_0/count[2]_net_1 ), .Y(
        \syn_md_module_1/syn_md_0/N_18 ));
    NOR2B \bri_dump_sw_0/reset_out_0  (.A(
        \bri_dump_sw_0/reset_out_5_net_1 ), .B(net_27), .Y(
        \bri_dump_sw_0/reset_out_0_net_1 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[7]_net_1 ));
    OR3 \scalestate_0/fst_lst_pulse_RNO_4  (.A(
        \scalestate_0/fst_lst_pulse8_NE_2 ), .B(
        \scalestate_0/fst_lst_pulse8_NE_1 ), .C(
        \scalestate_0/fst_lst_pulse8_NE_5 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_8 ));
    OR2A \scalestate_0/fst_lst_pulse_RNO  (.A(top_code_0_scale_rst_5), 
        .B(\scalestate_0/N_741 ), .Y(
        \scalestate_0/fst_lst_pulse_RNO_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[10]  (.A(
        \noisestate_0/acqtime[10]_net_1 ), .B(
        \noisestate_0/dectime[10]_net_1 ), .S(\noisestate_0/N_191 ), 
        .Y(\noisestate_0/N_67 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[5]  (.D(
        \DUMP_0/dump_coder_0/para2_4[5]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[5]_net_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[8]  (.A(
        \scanstate_0_timecount[8] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_246 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_54_i ));
    NOR3B \plusestate_0/timecount_1_RNO_1[3]  (.A(\plusestate_0/N_303 )
        , .B(top_code_0_pluse_rst_0), .C(\plusestate_0/CS[8]_net_1 ), 
        .Y(\plusestate_0/timecount_cnst[3] ));
    NOR2B \noisestate_0/rt_sw_RNO  (.A(\noisestate_0/N_110 ), .B(
        top_code_0_noise_rst), .Y(\noisestate_0/rt_sw_RNO_net_1 ));
    IOPAD_IN \ADC_pad[1]/U0/U0  (.PAD(ADC[1]), .Y(\ADC_pad[1]/U0/NET1 )
        );
    NOR2 \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[8]  (.A(
        \sd_acq_top_0/i_0[6] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[8]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_222 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/HND2_13_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net )
        , .C(\pd_pluse_top_0/count[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_13_net ));
    DFN1E1 \scanstate_0/dectime[1]  (.D(\top_code_0_scandata[1] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[1]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_71  (.D(
        \scalestate_0/timecount_20_iv_8[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[15] ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_1_inst  
        (.A(\pd_pluse_top_0/count_6[0] ), .B(
        \pd_pluse_top_0/count_6[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[1] ));
    OR3 \bridge_div_0/count_RNI3AD11[3]  (.A(
        \bridge_div_0/count[5]_net_1 ), .B(
        \bridge_div_0/count[4]_net_1 ), .C(
        \bridge_div_0/count[3]_net_1 ), .Y(
        \bridge_div_0/clear1_n17_NE_0[0] ));
    DFN1 \timer_top_0/timer_0/timedata[18]  (.D(
        \timer_top_0/timer_0/timedata_4[18] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[18]_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNICQ0I[7]  (.A(
        \sd_acq_top_0/count_3[7] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[7]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_22[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_5[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m187  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_186 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_187 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_188 ));
    DFN1E1 \scalestate_0/timecount_ret_10  (.D(
        \scalestate_0/timecount_cnst_m_0[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_cnst_m_0_reto[7] ));
    NOR2B \sd_acq_top_0/sd_sacq_state_0/cs_RNI1N9A[12]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[12]_net_1 ), .B(
        \sd_acq_top_0/i[9] ), .Y(\sd_acq_top_0/sd_sacq_state_0/N_230 ));
    DFN1 \scalestate_0/necount_LE_M  (.D(
        \scalestate_0/necount_LE_M_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount_LE_M_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m70_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[0] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i4_mux ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIAAC62[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_8[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_14[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_1[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_8[0] ));
    NOR3B \PLUSE_0/qq_coder_1/i_RNO[2]  (.A(bri_dump_sw_0_reset_out_0), 
        .B(\PLUSE_0/qq_coder_1/i_reg10_NE[0]_net_1 ), .C(
        \PLUSE_0/qq_coder_1/un1_qq_para2_i[0] ), .Y(
        \PLUSE_0/qq_coder_1/i_RNO_3[2] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_2_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ));
    NOR3B \top_code_0/k1_RNO_3  (.A(\top_code_0/N_13 ), .B(\xa_c[5] ), 
        .C(\top_code_0/N_158 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_5_i_a2_3 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[3]  (.D(
        \DUMP_0/dump_coder_0/para2_4[3]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[3]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[4]  (.A(
        \top_code_0_dumpdata_0[4] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[4]_net_1 ));
    DFN1 \topctrlchange_0/sw_acq2  (.D(\topctrlchange_0/sw_acq2_RNO_3 )
        , .CLK(GLA_net_1), .Q(sw_acq2_c));
    NOR2B \s_acq_change_0/s_acqnum_RNO[9]  (.A(\s_acq_change_0/N_79 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[9]_net_1 ));
    AO1C \plusestate_0/CS_RNO_0[4]  (.A(\plusestate_0/CS[3]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_srsts_i_0[4] ));
    NOR2 \top_code_0/un1_xa_8_16_i_i_o3_i_a2_3  (.A(\xa_c[13] ), .B(
        \xa_c[10] ), .Y(\top_code_0/un1_xa_8_16_i_i_o3_i_a2_3_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m104  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_101 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_104 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_105 ));
    DFN1E1 \scalestate_0/timecount_ret_59  (.D(
        \scalestate_0/timecount_20_iv_8[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[0] ));
    AOI1 \PLUSE_0/qq_state_1/cs_RNILLC8[4]  (.A(\PLUSE_0/i_2[3] ), .B(
        \PLUSE_0/qq_state_1/cs[3]_net_1 ), .C(
        \PLUSE_0/qq_state_1/cs[4]_net_1 ), .Y(
        \PLUSE_0/qq_state_1/N_84 ));
    IOBI_IB_OB_EB \xd_pad[14]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[14] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[14]/U0/NET3 ), .DOUT(
        \xd_pad[14]/U0/NET1 ), .EOUT(\xd_pad[14]/U0/NET2 ), .Y(
        \xd_in[14] ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_4  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_2_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_9_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_5_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_4_Y ));
    OR3 \top_code_0/scanload_RNO_0  (.A(\top_code_0/N_151 ), .B(
        \top_code_0/N_142 ), .C(\top_code_0/N_147 ), .Y(
        \top_code_0/N_202 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m6  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[1] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_7_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_62_i ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[0]  (.D(
        \top_code_0_state_1ms_data[0] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[0]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_69_RNO_0  (.A(
        \scalestate_0/CUTTIME180[15]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[15] ));
    MX2 \DSTimer_0/dump_sustain_timer_0/data_RNO_0[0]  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[0]_net_1 ), .B(
        \top_code_0_dump_sustain_data[0] ), .S(\DSTimer_0/AND2_0_Y ), 
        .Y(\DSTimer_0/dump_sustain_timer_0/N_24 ));
    OR3 \top_code_0/pluse_str_RNO_2  (.A(\top_code_0/N_328 ), .B(
        \top_code_0/N_327 ), .C(\top_code_0/N_319 ), .Y(
        \top_code_0/N_116 ));
    DFN1E1 \top_code_0/pd_pluse_data[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[10] ));
    NOR2B \top_code_0/pluse_str_RNO  (.A(\top_code_0/N_798 ), .B(
        net_27), .Y(\top_code_0/pluse_str_RNO_net_1 ));
    AO1A \scalestate_0/timecount_ret_2_RNO_2  (.A(
        \scalestate_0/N_1089 ), .B(\scalestate_0/S_DUMPTIME[6]_net_1 ), 
        .C(\scalestate_0/timecount_20_iv_1[6] ), .Y(
        \scalestate_0/timecount_20_iv_6[6] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[3]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_166  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_166_Y ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_68_i ));
    NOR3B \top_code_0/bri_datain_1_sqmuxa_0_a2  (.A(\top_code_0/N_331 )
        , .B(\top_code_0/N_332 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/bri_datain_1_sqmuxa ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[11]  (.A(
        \scalestate_0_timecount[11] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_198 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIUFK91[13]  (.A(
        \sd_acq_top_0/count_0[13] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[13]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_11[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_1[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[13]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[13]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_336 ));
    NOR3C \DUMP_0/dump_coder_0/i_RNO[4]  (.A(
        \DUMP_0/dump_coder_0/N_19 ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] ), .C(
        \DUMP_0/dump_coder_0/i_0_0_a2_0[4] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO[4]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m37  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_38_i ));
    NOR3 \DDS_0/dds_state_0/para_RNO[12]  (.A(
        \DDS_0/dds_state_0/N_333 ), .B(\DDS_0/dds_state_0/N_332 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[12] ), .Y(
        \DDS_0/dds_state_0/N_103 ));
    AO1C \state_1ms_0/timecount_RNO_3[6]  (.A(
        \state_1ms_0/M_DUMPTIME[6]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_i[0]_net_1 ), 
        .Y(\state_1ms_0/timecount_8_iv_0[6] ));
    MX2 \scan_scale_sw_0/s_start_RNO_0  (.A(
        \scan_scale_sw_0/s_start_5 ), .B(scan_scale_sw_0_s_start), .S(
        \top_code_0_change[1] ), .Y(\scan_scale_sw_0/N_26 ));
    AO1C \DUMP_0/dump_coder_0/un1_para114_5  (.A(
        \DUMP_0/dump_coder_0/para16_net_1 ), .B(
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ), .C(
        top_code_0_dumpload), .Y(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[0]_net_1 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[1]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[1] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[1]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_10  (.A(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[2]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m30  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_31 ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[5]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[5] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_1[5] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIV1ES[13]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[13]_net_1 ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_13[0] ));
    IOTRI_OB_EB \relay_close_pad[8]/U0/U1  (.D(\relay_close_c[8] ), .E(
        VCC), .DOUT(\relay_close_pad[8]/U0/NET1 ), .EOUT(
        \relay_close_pad[8]/U0/NET2 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[11]  (.D(
        \top_code_0_state_1ms_data[11] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[11]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m41_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[18] ));
    IOTRI_OB_EB \dumpon_pad/U0/U1  (.D(dumpon_c), .E(VCC), .DOUT(
        \dumpon_pad/U0/NET1 ), .EOUT(\dumpon_pad/U0/NET2 ));
    AO1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_59  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_60_i ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_0 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_8_0 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m46_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[13] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[13]  (.A(
        \state_1ms_0_timecount[13] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_192 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[5]  (.A(
        \top_code_0_dumpdata_0[5] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[5] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIUB452[4]  (.A(
        \ClockManagement_0/long_timer_0/count_c3 ), .B(
        \ClockManagement_0/long_timer_0/count[4]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c4 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m253  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[15] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_254 ));
    OR3 \scalestate_0/fst_lst_pulse_RNO_9  (.A(
        \scalestate_0/fst_lst_pulse8_0 ), .B(
        \scalestate_0/fst_lst_pulse8_2 ), .C(
        \scalestate_0/fst_lst_pulse8_9 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_5 ));
    DFN1E1 \top_code_0/pluseload  (.D(\top_code_0/N_90 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_pluseload));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[3] ));
    DFN1 \top_code_0/scale_rst_1_0  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_1));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m70  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m70_6 ));
    NOR2B \scalestate_0/timecount_20_iv_5_RNO_0[5]  (.A(
        \scalestate_0/OPENTIME_TEL[5]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[5] ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[0]  (.A(\s_acq_change_0/N_70 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[0]_net_1 ));
    NOR3A \PLUSE_0/bri_state_0/cs_RNO_0[2]  (.A(
        \PLUSE_0/bri_state_0/cs[0]_net_1 ), .B(\PLUSE_0/i_3[3] ), .C(
        \PLUSE_0/i_1[4] ), .Y(\PLUSE_0/bri_state_0/csse_1_0_a4_0_0 ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_16  (.A(
        \top_code_0_sigtimedata[13] ), .B(
        \ClockManagement_0/long_timer_0/count[13]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_13 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m14  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_13_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_14_0 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_15_0 ));
    NOR2 \PLUSE_0/bri_state_0/cs_RNO_7[3]  (.A(
        \PLUSE_0/bri_state_0/cs[3]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs[4]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_4 ));
    NOR3C \scalestate_0/S_DUMPTIME_1_sqmuxa_0_a2  (.A(
        \top_code_0_scalechoice_0_0[0] ), .B(\scalestate_0/N_60 ), .C(
        \scalestate_0/N_61 ), .Y(\scalestate_0/S_DUMPTIME_1_sqmuxa ));
    XOR2 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/UXOR2_12_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_15_net ), 
        .B(\pd_pluse_top_0/count[15] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[15] ));
    DFN1E1 \top_code_0/scaledatain[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[3] ));
    DFN1E1 \top_code_0/scalechoice[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/scalechoice_1_sqmuxa ), .Q(
        \top_code_0_scalechoice_0[0] ));
    DFN1E0 \DDS_0/dds_state_0/para[20]  (.D(\DDS_0/dds_state_0/N_123 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[20]_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI4N021[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_6[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIJAUE[0]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[0]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_0[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_100  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_100_Y ));
    DFN1E1 \top_code_0/noisedata[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[2] ));
    DFN1E1 \top_code_0/halfdata[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[3] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[2]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n2 ));
    DFN1E1 \top_code_0/change_0[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/change_1_sqmuxa ), .Q(
        \top_code_0_change_0[0] ));
    DFN1P0 \PLUSE_0/bri_state_0/cs[6]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_1[6] ), .CLK(ddsclkout_c), .PRE(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs_i_0[6] ));
    OR3 \scalestate_0/timecount_ret_23_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[10] ), .B(
        \scalestate_0/OPENTIME_TEL_m[10] ), .C(
        \scalestate_0/timecount_20_iv_4[10] ), .Y(
        \scalestate_0/timecount_20_iv_8[10] ));
    DFN1E1 \state_1ms_0/CUTTIME[19]  (.D(
        \top_code_0_state_1ms_data[3] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_380 ), .Q(\state_1ms_0/CUTTIME[19]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[4]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[9]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[9]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 )
        );
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m46 ));
    NOR3C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO_0[11]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c10 ));
    DFN1E1 \top_code_0/scandata[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[4] ));
    NOR3B \top_code_0/relay_on_1_sqmuxa_0_a2  (.A(\xa_c[6] ), .B(
        \top_code_0/relay_on_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_137 ), .Y(\top_code_0/relay_on_1_sqmuxa ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIGIDR2[9]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c8 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c10 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m145  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_146 ));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_23  (.A(
        \ClockManagement_0/clk_10k_0/count[0]_net_1 ), .B(
        \ClockManagement_0/clk_5M_en ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_partial_sum[0] ));
    AO1 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_44  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[1] )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[2] )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_COMP0_E[2] )
        );
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/PAND2_19_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), 
        .C(\sd_acq_top_0/count[16] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc1_25_net ));
    IOTRI_OB_EB \GLA_pad/U0/U1  (.D(GLA_net_1), .E(VCC), .DOUT(
        \GLA_pad/U0/NET1 ), .EOUT(\GLA_pad/U0/NET2 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIUJCM[3]  (.A(
        \sd_acq_top_0/count_10[3] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[3]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_0_0[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_10[0] ));
    IOPAD_TRI \relay_on_pad[2]/U0/U0  (.D(\relay_on_pad[2]/U0/NET1 ), 
        .E(\relay_on_pad[2]/U0/NET2 ), .PAD(relay_on[2]));
    DFN1E0 \DUMP_0/dump_coder_0/para4[2]  (.D(
        \DUMP_0/dump_coder_0/para4_4[2]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[2]_net_1 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[6]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c4 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n6 ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[0] ), .CLK(
        GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ));
    DFN1 \scalestate_0/s_acqnum_1[10]  (.D(
        \scalestate_0/s_acqnum_1_RNO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[10] ));
    DFN1E1 \top_code_0/state_1ms_data[5]  (.D(\GPMI_0_dataout[5] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[5] ));
    NOR2A \scalestate_0/timecount_ret_28_RNO_0  (.A(
        \scalestate_0/S_DUMPTIME[1]_net_1 ), .B(\scalestate_0/N_1089 ), 
        .Y(\scalestate_0/S_DUMPTIME_m[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m184  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_183 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_184 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_185 ));
    DFN1E1 \scanstate_0/dectime[3]  (.D(\top_code_0_scandata[3] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[3]_net_1 ));
    NOR2A \top_code_0/pn_change_RNO_1  (.A(\top_code_0/N_340 ), .B(
        \top_code_0/N_148 ), .Y(\top_code_0/N_300 ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_i[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_21[10] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO[10]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[12]_net_1 )
        );
    OA1C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[6]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/en2 ), .B(
        \pd_pluse_top_0/i_0[4] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs[5]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_186 ));
    IOPAD_IN \xa_pad[11]/U0/U0  (.PAD(xa[11]), .Y(\xa_pad[11]/U0/NET1 )
        );
    OR3 \timer_top_0/state_switch_0/dataout_RNO[12]  (.A(
        \timer_top_0/state_switch_0/N_255 ), .B(
        \timer_top_0/state_switch_0/N_256 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[12] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[12]_net_1 ));
    AO1A \scalestate_0/timecount_ret_73_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[7]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[7] ), .Y(
        \scalestate_0/timecount_20_iv_0[7] ));
    NOR3 \top_code_0/inv_turn_RNO_2  (.A(\top_code_0/N_144 ), .B(
        \top_code_0/N_167 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/N_322 ));
    NOR2B \state_1ms_0/dump_start_RNO  (.A(\state_1ms_0/N_87 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/dump_start_RNO_2_net_1 ));
    MX2 \nsctrl_choice_0/sw_acq2_RNO_0  (.A(scanstate_0_sw_acq2), .B(
        noisestate_0_sw_acq2), .S(top_code_0_n_s_ctrl_0), .Y(
        \nsctrl_choice_0/sw_acq2_5 ));
    NOR2 \plusestate_0/CS_RNIDNHP[1]  (.A(\plusestate_0/CS[2]_net_1 ), 
        .B(\plusestate_0/CS[1]_net_1 ), .Y(\plusestate_0/N_303 ));
    NOR3C \DUMP_ON_0/off_on_state_0/cs_RNO[0]  (.A(
        \DUMP_ON_0/off_on_state_0/N_42_i ), .B(\DUMP_ON_0/i_5[0] ), .C(
        OR2_2_Y), .Y(\DUMP_ON_0/off_on_state_0/N_36_i ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_54  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[9] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[12] ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[13] ));
    NOR2A \PLUSE_0/bri_state_0/cs_RNO_0[11]  (.A(
        \PLUSE_0/bri_state_0/cs[10]_net_1 ), .B(
        \PLUSE_0/bri_state_0/N_142 ), .Y(
        \PLUSE_0/bri_state_0/csse_10_0_a4_0_0 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[9]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c8 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n9 ));
    NOR3C \scalestate_0/timecount_ret_14_RNO_1  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[9]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[9] ));
    DFN1E1 \plusestate_0/timecount_1[15]  (.D(
        \plusestate_0/timecount_5[15] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[15] ));
    NOR3A \topctrlchange_0/rt_sw_RNO_2  (.A(nsctrl_choice_0_rt_sw), .B(
        \top_code_0_change_0[0] ), .C(\top_code_0_change[1] ), .Y(
        \topctrlchange_0/rt_swin1_m ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/ADD_20x20_slow_I19_Y )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[19] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[9]  (.D(
        \top_code_0_sd_sacq_data[9] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[9]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[2]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[12]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[12]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[12] ));
    DFN1 \DUMP_ON_0/off_on_timer_0/count[3]  (.D(
        \DUMP_ON_0/off_on_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/count_5[3] ));
    MX2 \scalestate_0/CS_RNO_0[10]  (.A(\scalestate_0/CS[10]_net_1 ), 
        .B(\scalestate_0/CS[20]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1224 ));
    NOR2B \DUMP_0/off_on_timer_1/count_RNIEPL21[2]  (.A(
        \DUMP_0/off_on_timer_1/count_c1 ), .B(\DUMP_0/count_0[2] ), .Y(
        \DUMP_0/off_on_timer_1/count_c2 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[6]  (.D(
        \top_code_0_state_1ms_data[6] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[6]_net_1 ));
    DFN1E1 \noisestate_0/dectime[14]  (.D(\top_code_0_noisedata[14] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[14]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIRVS7[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[1]_net_1 ), .B(
        \sd_acq_top_0/count_10[1] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_1[0] ));
    DFN1E1 \scalestate_0/timecount_ret_63  (.D(
        \scalestate_0/timecount_20_iv_7[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[13] ));
    NOR2B \topctrlchange_0/interupt_RNO_3  (.A(
        plusestate_0_state_over_n), .B(\top_code_0_change[1] ), .Y(
        \topctrlchange_0/interin3_m ));
    DFN1E1 \scalestate_0/S_DUMPTIME[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[10]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIOTC81[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c2 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c4 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m38  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_37 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_38 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_39 ));
    DFN1E0 \DDS_0/dds_state_0/para[19]  (.D(\DDS_0/dds_state_0/N_165 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[19]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_2_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_122_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_118_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_2_inst ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_9_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_11_net ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[11] ));
    DFN1 \DUMP_0/off_on_timer_1/count[2]  (.D(
        \DUMP_0/off_on_timer_1/count_n2 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[2] ));
    NOR2A \DDS_0/dds_coder_0/m3_e_1  (.A(dds_change_0_dds_rst), .B(
        \DDS_0/count[0] ), .Y(\DDS_0/dds_coder_0/m3_e_1_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_RNO_0  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_entop ), 
        .B(scan_scale_sw_0_s_start), .C(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/clkout_1_sqmuxa )
        );
    DFN1E1 \scalestate_0/PLUSETIME180[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[14]_net_1 ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[1]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_33_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[1] ));
    NOR2B \scalestate_0/timecount_ret_81_RNO_0  (.A(
        \scalestate_0/OPENTIME[4]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[4] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[2]  (.A(
        \noisestate_0_timecount[2] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_230 ));
    NOR2B \scalestate_0/timecount_ret_73_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[7]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[7] ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[6]  (.A(
        \DUMP_0/dump_timer_0/count_c5 ), .B(\DUMP_0/count_0[6] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n6 ));
    AX1C \timer_top_0/timer_0/un2_timedata_I_12  (.A(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .C(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .Y(
        \timer_top_0/timer_0/I_12_2 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_56_i ));
    DFN1E1 \top_code_0/scaledatain[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[0] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_39_i ));
    DFN1E1 \scalestate_0/CUTTIMEI90[19]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[19]_net_1 )
        );
    NOR2A \DUMP_0/dump_coder_0/para4_4[9]  (.A(
        \top_code_0_dumpdata_0[9] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[9]_net_1 ));
    DFN1 \PLUSE_0/qq_timer_0/count[0]  (.D(
        \PLUSE_0/qq_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_9[0] ));
    NOR3B \top_code_0/scalechoice_1_sqmuxa_0_a2  (.A(
        \top_code_0/N_331 ), .B(\top_code_0/N_332 ), .C(
        \top_code_0/N_165 ), .Y(\top_code_0/scalechoice_1_sqmuxa ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[3]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[2] ), 
        .Y(\DDS_0/dds_state_0/N_489 ));
    OR3 \scalestate_0/timecount_ret_2_RNO  (.A(
        \scalestate_0/timecount_20_iv_3[6] ), .B(
        \scalestate_0/timecount_20_iv_2[6] ), .C(
        \scalestate_0/timecount_20_iv_6[6] ), .Y(
        \scalestate_0/timecount_20_iv_9[6] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[2]_net_1 ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[2]  (.A(
        \DUMP_0/dump_timer_0/count_c1 ), .B(\DUMP_0/count_1[2] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n2 ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNIB0MS[11]  (.A(
        \DUMP_0/dump_coder_0/para2[11]_net_1 ), .B(\DUMP_0/count[11] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_11[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[1]  (.A(
        \state_1ms_0_timecount[1] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_237 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_66_i ));
    AO1 \scalestate_0/necount_cmp_0/AO1_1  (.A(
        \scalestate_0/necount_cmp_0/AND3_2_Y ), .B(
        \scalestate_0/necount_cmp_0/NAND3A_4_Y ), .C(
        \scalestate_0/necount_cmp_0/NAND3A_0_Y ), .Y(
        \scalestate_0/necount_cmp_0/AO1_1_Y ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[4]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[4] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[15]_net_1 )
        );
    DFN1E1 \state_1ms_0/PLUSETIME[4]  (.D(
        \top_code_0_state_1ms_data[4] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[4]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m166  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_167 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[10]  (.A(
        \s_acq_change_0/s_acqnum_5[10] ), .B(
        \s_acq_change_0_s_acqnum[10] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_80 ));
    DFN1E1 \plusestate_0/DUMPTIME[11]  (.D(\top_code_0_plusedata[11] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[11]_net_1 ));
    DFN1E1 \top_code_0/s_addchoice[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice[0] ));
    OR3 \state_1ms_0/timecount_RNO_1[14]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[14] ), .B(
        \state_1ms_0/CUTTIME_m[14] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[14] ), .Y(
        \state_1ms_0/timecount_8[14] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[2]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[3]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_488 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[10]  (.A(
        \ClockManagement_0/long_timer_0/count_c9 ), .B(
        \ClockManagement_0/long_timer_0/count[10]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n10 ));
    NOR2 \syn_md_module_1/syn_md_0/syn_md_out_RNO_0  (.A(syn_md_out_c), 
        .B(\syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en ), .Y(
        \syn_md_module_1/syn_md_0/N_30 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[9]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_54_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[9] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[11]  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c10 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n11 ));
    NOR2B \state_1ms_0/timecount_RNO_6[1]  (.A(
        \state_1ms_0/CUTTIME[1]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[1] ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[2]  (.A(s_acq180_c), .B(
        net_27), .Y(\sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[2] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m276  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_277 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_60  (.A(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[15] ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIINCT3[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_2 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_1 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_7 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_11 )
        );
    NOR3B \top_code_0/un1_state_1ms_rst_n117_i_a2  (.A(\xa_c[7] ), .B(
        \top_code_0/un1_state_1ms_rst_n117_i_a2_0_net_1 ), .C(
        \top_code_0/N_139 ), .Y(\top_code_0/N_264 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[5]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[6]  (.D(
        \DUMP_0/dump_coder_0/para4_4[6]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[6]_net_1 ));
    MX2 \scanstate_0/timecount_1_RNO_0[8]  (.A(
        \scanstate_0/acqtime[8]_net_1 ), .B(
        \scanstate_0/dectime[8]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_66 ));
    XA1A \scalestate_0/necount_cmp_0/AND2_0  (.A(
        \scalestate_0/M_NUM[10]_net_1 ), .B(
        \scalestate_0/necount[10]_net_1 ), .C(
        \scalestate_0/necount_cmp_0/XNOR2_2_Y ), .Y(
        \scalestate_0/necount_cmp_0/AND2_0_Y ));
    NOR3B \scalestate_0/CS_RNI4LFN[12]  (.A(
        \scalestate_0/CS[12]_net_1 ), .B(top_code_0_scale_rst_1), .C(
        scalestate_0_ne_le), .Y(\scalestate_0/N_252 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[7]  (.D(
        \DUMP_0/dump_coder_0/para4_4[7]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[7]_net_1 ));
    OR3A \top_code_0/pluse_lc_3_i_o2  (.A(\xa_c[7] ), .B(
        \top_code_0/N_139 ), .C(\top_code_0/N_144 ), .Y(
        \top_code_0/N_175 ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/fAND2_8_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_2_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ), 
        .C(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_10_net )
        , .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_9_net ));
    NOR3 \top_code_0/dumpload_RNO_1  (.A(\top_code_0/N_144 ), .B(
        \top_code_0/N_148 ), .C(\top_code_0/N_165 ), .Y(
        \top_code_0/N_278 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[6]  (.A(\s_acq_change_0/N_76 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[6]_net_1 ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n3 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        );
    MX2 \scanstate_0/timecount_1_RNO[8]  (.A(\scanstate_0/N_66 ), .B(
        \scanstate_0/timecount_cnst[4] ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[8] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[5]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[4] ), 
        .Y(\DDS_0/dds_state_0/N_319 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_161  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_155_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_115_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_161_Y ));
    AO1 \bridge_div_0/dataall_1_I_16  (.A(
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0_1[0] ), .B(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_1[0] ), .C(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_2[0] ), .Y(
        \bridge_div_0/dataall_1[3] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[2]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n2 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[9]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n9 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ));
    AO1B \noisestate_0/CS_RNO_0[1]  (.A(\noisestate_0/CS_li[0] ), .B(
        timer_top_0_clk_en_noise), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/CS_srsts_i_0[1] ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_10  
        (.A(\s_acq_change_0_s_stripnum[0] ), .B(
        \s_acq_change_0_s_stripnum[1] ), .C(
        \s_acq_change_0_s_stripnum[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[0] )
        );
    IOPAD_IN \xa_pad[12]/U0/U0  (.PAD(xa[12]), .Y(\xa_pad[12]/U0/NET1 )
        );
    AND3B \sd_acq_top_0/sd_sacq_state_0/cs_RNIDTT7[11]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[4]_net_1 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[11]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/ns_0_1_i_a2_0 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_245 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_5_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_140_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_48_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_5_inst ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_2_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_2_net ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[0]_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[17]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[17] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[17] ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_1  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_0_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_6_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_3_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_1_Y ));
    OR3 \state_1ms_0/timecount_RNO_1[12]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[12] ), .B(
        \state_1ms_0/CUTTIME_m[12] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[12] ), .Y(
        \state_1ms_0/timecount_8[12] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[23]  (.D(
        \top_code_0_dds_configdata[6] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[23]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_choice[3]  (.D(\GPMI_0_dataout[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_choice_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_choice[3] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[6]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c4 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n6 ));
    DFN1 \scanstate_0/CS[1]  (.D(\scanstate_0/CS_RNO_2[1] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[1]_net_1 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNICI142[7]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_11[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_13[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_13[0] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[0]  (.A(
        \scalestate_0_strippluse[0] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m292  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_291 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_292 ), .S(
        \top_code_0_s_addchoice[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_293 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[6]  (.D(
        \ClockManagement_0/long_timer_0/count_n6 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[6]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[1]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        , .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m79  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_80 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[7]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_20_0 ), .Y(
        \timer_top_0/timer_0/timedata_4[7] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m120  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[19] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_121 ));
    NOR2 \DUMP_0/off_on_coder_1/i_RNO_1[1]  (.A(\DUMP_0/count_2[0] ), 
        .B(\DUMP_0/count_2[1] ), .Y(\DUMP_0/off_on_coder_1/i_0_1[1] ));
    NOR2A \state_1ms_0/timecount_RNO_6[6]  (.A(
        \state_1ms_0/CS[8]_net_1 ), .B(\state_1ms_0/CUTTIME[6]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_i_m[6] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m178  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_179 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[7]  (.D(
        \DUMP_0/dump_coder_0/para2_4[7]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[7]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m70_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[0] ));
    OR3 \scalestate_0/timecount_ret_28_RNI70O  (.A(
        \scalestate_0/timecount_20_iv_9_reto[1] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[1] ), .C(
        \scalestate_0/timecount_cnst_m_reto[1] ), .Y(
        \scalestate_0_timecount[1] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[8]  (.D(
        \top_code_0_pd_pluse_data[8] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[8]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[28]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[29]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_480 ));
    DFN1E1 \top_code_0/bri_datain[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[0] ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[3]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIJUOK[4]  (.A(
        \DUMP_0/dump_coder_0/para6[4]_net_1 ), .B(\DUMP_0/count_1[4] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_4[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m45_4 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[14] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/ADD_20x20_slow_I19_Y_5 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[19] ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_100_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_1_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ));
    DFN1E1 \scalestate_0/timecount_ret_56  (.D(
        \scalestate_0/timecount_20_0_iv_4[19] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_4_reto[19] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[1]  (.D(
        \top_code_0_pd_pluse_data[1] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[1]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m43_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] ));
    XA1 \PLUSE_0/qq_timer_1/count_RNO[1]  (.A(\PLUSE_0/count_7[1] ), 
        .B(\PLUSE_0/count_7[0] ), .C(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_1/count_n1 ));
    DFN1E1 \top_code_0/sd_sacq_choice[1]  (.D(\GPMI_0_dataout[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_choice_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_choice[1] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[9]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c8 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n9 ));
    XOR2 \scalestate_0/M_pulse_RNO_10  (.A(
        \scalestate_0/M_NUM[1]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .Y(\scalestate_0/M_pulse8_1 )
        );
    IOPAD_BI \xd_pad[15]/U0/U0  (.D(\xd_pad[15]/U0/NET1 ), .E(
        \xd_pad[15]/U0/NET2 ), .Y(\xd_pad[15]/U0/NET3 ), .PAD(xd[15]));
    DFN1 \top_code_0/state_1ms_rst_n  (.D(
        \top_code_0/state_1ms_rst_n_0_0_RNI848T5_net_1 ), .CLK(
        GLA_net_1), .Q(top_code_0_state_1ms_rst_n));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_70_i ));
    AO1 \state_1ms_0/timecount_RNO_2[10]  (.A(
        \state_1ms_0/M_DUMPTIME[10]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[10] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[10] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_18  (.A(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[5]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[5]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_66_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[14]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[14] ));
    NOR2A \scalestate_0/strippluse_RNO_1[0]  (.A(\scalestate_0/N_420 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[0] ));
    NOR2B \scalestate_0/timecount_ret_20_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[8]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[8] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[20]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[21]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_468 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIMQ9N1[3]  (.A(
        \ClockManagement_0/long_timer_0/count_c2 ), .B(
        \ClockManagement_0/long_timer_0/count[3]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c3 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_2  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_1_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_1_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_3_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_2_Y ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[0]  (.A(
        \scalestate_0/s_acqnum_7[0] ), .B(\scalestate_0_s_acqnum[0] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_547 ));
    DFN1 \scalestate_0/s_acqnum_1[2]  (.D(
        \scalestate_0/s_acqnum_1_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[2] ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/M_NUM[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_3_Y ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[25]  (.A(
        \top_code_0_dds_configdata[8] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_307 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[25] ));
    DFN1 \ClockManagement_0/clk_10k_0/clock_10khz  (.D(
        \ClockManagement_0/clk_10k_0/clock_10khz_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(clock_10khz));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[3]_net_1 ));
    OR2 \PLUSE_0/bri_coder_0/un2lto7_1  (.A(\PLUSE_0/count_2[6] ), .B(
        \PLUSE_0/count_8[3] ), .Y(
        \PLUSE_0/bri_coder_0/un2lto7_1_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_state_0/cs_RNO[4]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/en1 ), .B(\sd_acq_top_0/i_1[5] ), 
        .C(\sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_5[4] ));
    NOR2B \scalestate_0/CS_RNO[20]  (.A(\scalestate_0/N_1232 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/CS_RNO[20]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_0  (.A(\ADC_c[10] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[29]  (.A(
        \top_code_0_dds_configdata[12] ), .B(\DDS_0/dds_state_0/N_569 )
        , .C(\DDS_0/dds_state_0/N_482 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[29] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[25]  (.A(
        \DDS_0/dds_state_0/N_310 ), .B(\DDS_0/dds_state_0/N_309 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[25] ), .Y(
        \DDS_0/dds_state_0/N_25 ));
    DFN1 \CAL_0/cal_div_0/count[3]  (.D(\CAL_0/cal_div_0/count_5[3] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[3]_net_1 ));
    XO1 \DUMP_0/dump_coder_0/para2_RNIKQO01[2]  (.A(
        \DUMP_0/count_1[2] ), .B(\DUMP_0/dump_coder_0/para2[2]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_3_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_3[0] ));
    IOIN_IB \xa_pad[0]/U0/U1  (.YIN(\xa_pad[0]/U0/NET1 ), .Y(\xa_c[0] )
        );
    NOR3B \scalestate_0/OPENTIME_452_e  (.A(\scalestate_0/N_62 ), .B(
        \scalestate_0/N_65 ), .C(\top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/N_1665 ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_5  (.A(
        \scalestate_0/necount[7]_net_1 ), .B(
        \scalestate_0/M_NUM[7]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_5_Y ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[6]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[6] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n7 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7]/Y ));
    NOR3C \ClockManagement_0/long_timer_0/timeup_RNO_3  (.A(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_2 ), .B(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_1 ), .C(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_10 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_13 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[10]_net_1 ));
    DFN1E1 \scalestate_0/PLUSETIME180[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[0]_net_1 ));
    DFN1E1 \scanstate_0/dectime[14]  (.D(\top_code_0_scandata[14] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[14]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i10_mux ));
    XOR2 \ClockManagement_0/long_timer_0/timeup_RNO_9  (.A(
        \top_code_0_sigtimedata[9] ), .B(
        \ClockManagement_0/long_timer_0/count[9]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clear_n4_9 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_6_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_66_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_77_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_9_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_6_inst ));
    AO1A \scalestate_0/timecount_ret_59_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[0]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[0] ), .Y(
        \scalestate_0/timecount_20_iv_0[0] ));
    AOI1 \DUMP_ON_0/off_on_state_0/cs_RNI413F[1]  (.A(
        DUMP_ON_0_dump_on), .B(\DUMP_ON_0/i_5[1] ), .C(
        \DUMP_ON_0/off_on_state_0/cs[1]_net_1 ), .Y(
        \DUMP_ON_0/off_on_state_0/N_42_i ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_11  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[8] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/N_2 ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIKD1G[0]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[0]_net_1 ), 
        .B(\pd_pluse_top_0/count_6[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_0[0] ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_62  (.A(
        \timer_top_0/timer_0/N_2 ), .B(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .Y(
        \timer_top_0/timer_0/I_62 ));
    DFN1 \DUMP_OFF_0/off_on_coder_0/i[0]  (.D(
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/i_3[0] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m70  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m70_5 ));
    OR3 \scalestate_0/M_pulse_RNO_9  (.A(\scalestate_0/M_pulse8_0 ), 
        .B(\scalestate_0/M_pulse8_2 ), .C(\scalestate_0/M_pulse8_9 ), 
        .Y(\scalestate_0/M_pulse8_NE_5 ));
    AX1C \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/POR2_9_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), .C(
        \sd_acq_top_0/count_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[12] ));
    DFN1E1 \top_code_0/sd_sacq_data[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[10] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_68_i ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_144  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_144_Y ));
    OR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_2  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[2]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_3_0 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNISD6K[3]  (.A(
        \sd_acq_top_0/count_10[3] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[3]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_0_0[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_10[0] ));
    DFN1E1 \top_code_0/RAM_Rd_rst  (.D(\top_code_0/N_58 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_RAM_Rd_rst));
    AO1C \state_1ms_0/timecount_RNO_3[2]  (.A(
        \state_1ms_0/M_DUMPTIME[2]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_i[0]_net_1 ), 
        .Y(\state_1ms_0/timecount_8_iv_0[2] ));
    NOR2A \PLUSE_0/qq_state_0/cs_RNO[4]  (.A(\PLUSE_0/qq_state_0/cs4 ), 
        .B(\PLUSE_0/qq_state_0/N_84 ), .Y(
        \PLUSE_0/qq_state_0/cs_RNO_2[4] ));
    XA1 \DUMP_0/off_on_timer_0/count_RNO[2]  (.A(\DUMP_0/count_2[2] ), 
        .B(\DUMP_0/off_on_timer_0/count_c1 ), .C(
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_0/count_n2 ));
    NOR2B \scalestate_0/pn_out_RNO  (.A(\scalestate_0/N_571 ), .B(
        top_code_0_scale_rst), .Y(\scalestate_0/pn_out_RNO_net_1 ));
    DFN1P0 \PLUSE_0/bri_state_0/cs[7]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_0[7] ), .CLK(ddsclkout_c), .PRE(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs_i_0[7] ));
    DFN1E1 \top_code_0/state_1ms_data[8]  (.D(\GPMI_0_dataout[8] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[8] ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[4]  (.D(
        \top_code_0_cal_data[4] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[4] ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/PXOR2_13_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_17_net ), 
        .B(\sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[17] ));
    DFN1E1 \top_code_0/dds_configdata[0]  (.D(\GPMI_0_dataout[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[0] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_56_i ));
    DFN1E1 \scalestate_0/DUMPTIME[8]  (.D(\top_code_0_scaledatain[8] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[8]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[1]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[1] ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_3  (.A(
        \scalestate_0/M_NUM[7]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .C(
        \scalestate_0/necount_cmp_0/OR2A_2_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_3_Y ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI04P21[12]  (.A(
        \sd_acq_top_0/count_0[12] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[12]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_7[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[21]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[21]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_510 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[5]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[10]  (.A(
        \state_1ms_0/PLUSECYCLE[10]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[10] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_75  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_75_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_79  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_79_Y ));
    DFN1 \scalestate_0/CS_0[11]  (.D(
        \scalestate_0/CS_RNIRUEO[10]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/CS_0[11]_net_1 ));
    MX2 \top_code_0/relay_close_RNO_0[1]  (.A(\relay_close_c[1] ), .B(
        \GPMI_0_dataout_0[1] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_820 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[15]  (.A(
        \noisestate_0_timecount[15] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_185 ));
    DFN1E1 \plusestate_0/PLUSETIME[13]  (.D(\top_code_0_plusedata[13] )
        , .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[13]_net_1 ));
    DFN1E1 \top_code_0/s_addchoice_4[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_4[0] ));
    DFN1 \scalestate_0/load_out  (.D(\scalestate_0/load_out_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(scalestate_0_load_out));
    DFN1E1 \noisestate_0/acqtime[13]  (.D(\top_code_0_noisedata[13] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[13]_net_1 ));
    NOR3C \DUMP_0/off_on_state_1/cs_RNO[0]  (.A(
        state1ms_choice_0_reset_out), .B(\DUMP_0/i_0[0] ), .C(
        \DUMP_0/off_on_state_1/N_42_i ), .Y(
        \DUMP_0/off_on_state_1/N_36_i ));
    AO1C \DUMP_0/dump_coder_0/un1_para114_2  (.A(
        \DUMP_0/dump_coder_0/para19_net_1 ), .B(
        \DUMP_0/dump_coder_0/un1_dump_choice_2_net_1 ), .C(
        top_code_0_dumpload), .Y(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_39  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[8] ), .Y(
        \timer_top_0/timer_0/N_9 ));
    MX2 \noisestate_0/timecount_1_RNO_0[7]  (.A(
        \noisestate_0/acqtime[7]_net_1 ), .B(
        \noisestate_0/dectime[7]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_64 ));
    RAM512X18 #( .MEMORYFILE("RAM_R7C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R7C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_7_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_7_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_0_net ));
    DFN1E1 \scanstate_0/timecount_1[6]  (.D(
        \scanstate_0/timecount_5[6] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[6] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[17]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[17]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m7  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i2_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[2] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i4_mux ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI4MCH[13]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[13]_net_1 ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_13[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[26]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[27]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_472 ));
    NOR3C \scalestate_0/timecount_ret_1_RNO_3  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[5]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[5] ));
    AO1 \scalestate_0/timecount_ret_63_RNO_2  (.A(
        \scalestate_0/CUTTIME180_TEL[13]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[13] )
        , .Y(\scalestate_0/timecount_20_iv_3[13] ));
    DFN1E1 \scanstate_0/timecount_1[2]  (.D(
        \scanstate_0/timecount_5[2] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[2] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[5]  (.A(
        \timer_top_0/state_switch_0/N_217 ), .B(
        \timer_top_0/state_switch_0/N_219 ), .C(
        \timer_top_0/state_switch_0/N_218 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[5] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m246  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_247 ));
    NOR3C \PLUSE_0/bri_state_0/cs_RNO_4[3]  (.A(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_4 ), .B(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_3 ), .C(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_7 ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_10 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[0]  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_e0 ));
    DFN1E1 \top_code_0/n_s_ctrl  (.D(\top_code_0/N_76 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_n_s_ctrl));
    DFN1 \timer_top_0/timer_0/timedata[15]  (.D(
        \timer_top_0/timer_0/timedata_4[15] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[15]_net_1 ));
    IOTRI_OR_EB \ddsdata_pad/U0/U1  (.D(\DDS_0/dds_state_0/N_21 ), .E(
        VCC), .OCLK(GLA_net_1), .DOUT(\ddsdata_pad/U0/NET1 ), .EOUT(
        \ddsdata_pad/U0/NET2 ));
    DFN1E1 \state_1ms_0/CUTTIME[16]  (.D(
        \top_code_0_state_1ms_data[0] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_380 ), .Q(\state_1ms_0/CUTTIME[16]_net_1 ));
    NOR2B \bri_dump_sw_0/phase_ctr_RNO  (.A(
        \bri_dump_sw_0/phase_ctr_5 ), .B(net_27), .Y(
        \bri_dump_sw_0/phase_ctr_RNO_net_1 ));
    DFN1E1 \top_code_0/n_acqnum[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_87  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_124_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_2_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_87_Y ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[9]  (.A(
        \DDS_0/dds_state_0/para[9]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_286 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[9] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_9  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_119_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_57_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_9_Y ));
    IOIN_IB \ADC_pad[4]/U0/U1  (.YIN(\ADC_pad[4]/U0/NET1 ), .Y(
        \ADC_c[4] ));
    AO1 \scalestate_0/timecount_ret_54_RNO  (.A(
        \scalestate_0/OPENTIME[19]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[19] ), .Y(
        \scalestate_0/timecount_20_0_iv_0[19] ));
    DFN1E1 \top_code_0/plusedata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[7] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[7]  (.A(
        \timer_top_0/state_switch_0/N_207 ), .B(
        \timer_top_0/state_switch_0/N_209 ), .C(
        \timer_top_0/state_switch_0/N_208 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[7] ));
    MX2 \scanstate_0/timecount_1_RNO[5]  (.A(\scanstate_0/N_63 ), .B(
        net_33_0), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[5] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m16  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_17_0 ));
    XA1 \DUMP_ON_0/off_on_timer_0/count_RNO[1]  (.A(
        \DUMP_ON_0/count_5[1] ), .B(\DUMP_ON_0/count_5[0] ), .C(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_n1 ));
    OA1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_58  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_58_i ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_3_0 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_7_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_68_i ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[5] ));
    AND2A \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y ));
    DFN1 \top_code_0/pluse_rst  (.D(
        \top_code_0/pluse_rst_0_0_RNIO7ND3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_pluse_rst));
    NOR3C \scalestate_0/timecount_ret_73_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[7]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[7] ));
    OR2 \scalestate_0/timecount_20_iv_8[4]  (.A(
        \scalestate_0/timecount_20_iv_5[4]_net_1 ), .B(
        \scalestate_0/timecount_20_iv_4[4]_net_1 ), .Y(
        \scalestate_0/timecount_20_iv_8[4]_net_1 ));
    DFN1 \state_1ms_0/timecount[17]  (.D(
        \state_1ms_0/timecount_RNO[17]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[17] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_90  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_90_Y ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/TND2_15_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_22_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_15_net ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[14]_net_1 ));
    OA1B \scanstate_0/CS_RNO[5]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[5]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[5] ), 
        .Y(\scanstate_0/CS_RNO_2[5] ));
    MX2 \plusestate_0/timecount_1_RNO_0[4]  (.A(
        \plusestate_0/PLUSETIME[4]_net_1 ), .B(
        \plusestate_0/DUMPTIME[4]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_75 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[2]_net_1 ));
    DFN1 \DDS_0/dds_state_0/state_over  (.D(
        \DDS_0/dds_state_0/state_over_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0_state_over ));
    IOPAD_IN \xa_pad[14]/U0/U0  (.PAD(xa[14]), .Y(\xa_pad[14]/U0/NET1 )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_82  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_82_Y ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI4F6B[4]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_4[0] ));
    IOIN_IB \ADC_pad[8]/U0/U1  (.YIN(\ADC_pad[8]/U0/NET1 ), .Y(
        \ADC_c[8] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_102  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_13_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_71_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_102_Y ));
    NOR3C \DUMP_OFF_0/off_on_state_0/cs_RNO[0]  (.A(
        \DUMP_OFF_0/off_on_state_0/N_42_i ), .B(\DUMP_OFF_0/i_3[0] ), 
        .C(bri_dump_sw_0_reset_out_0), .Y(
        \DUMP_OFF_0/off_on_state_0/N_36_i ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[12]  (.A(
        \noisestate_0_timecount[12] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_255 ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[11]  (.A(
        \PLUSE_0/bri_state_0/cs[11]_net_1 ), .B(
        \PLUSE_0/bri_state_0/csse_10_0_a4_0_0 ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[11] ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m22  
        (.A(\s_acq_change_0_s_stripnum[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[7]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i14_mux )
        );
    DFN1E1 \scalestate_0/timecount_ret_17  (.D(
        \scalestate_0/un1_timecount_2_sqmuxa_1 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/un1_timecount_2_sqmuxa_1_reto ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[21]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1789 ), .Q(
        \scalestate_0/OPENTIME_TEL[21]_net_1 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[1]  (.D(
        \PLUSE_0/bri_state_0/cs_ns_e[1] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[1]_net_1 ));
    OR2 \top_code_0/scaleload_RNO_0  (.A(\top_code_0/N_174 ), .B(
        \top_code_0/N_147 ), .Y(\top_code_0/N_217 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m228  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_229 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m165  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_162 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_165 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_166 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI2M063[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_5[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_4[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_11[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_13[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[8]  (.D(
        \DUMP_0/dump_coder_0/para5_4[8] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[8]_net_1 ));
    NOR3B \scalestate_0/CUTTIME180_TEL_494_e  (.A(\scalestate_0/N_61 ), 
        .B(\scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 ), .C(
        \top_code_0_scalechoice_0_0[0] ), .Y(\scalestate_0/N_1707 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m13  
        (.A(\s_acq_change_0_s_stripnum[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[4]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i8_mux ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_ADD_16x16_slow_I15_Y  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[14]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_37_i ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[15]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y )
        );
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_6  (.A(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .B(
        \timer_top_0/dataout[19] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_6_Y ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[3]  (.A(
        \scalestate_0_strippluse[3] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[3] ));
    DFN1E1 \scalestate_0/PLUSETIME180[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[3]_net_1 ));
    NOR2B \ClockManagement_0/clk_10k_0/clock_10khz_RNO  (.A(net_27), 
        .B(\ClockManagement_0/clk_10k_0/clock_10khz_RNO_0_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/clock_10khz_RNO_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_81  (.D(
        \scalestate_0/timecount_20_iv_2[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_2_reto[4] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m148  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_149 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[15]_net_1 ));
    DFN1 \scalestate_0/necount[7]  (.D(
        \scalestate_0/necount_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[7]_net_1 ));
    MX2 \state_1ms_0/rt_sw_RNO_0  (.A(state_1ms_0_rt_sw), .B(
        \state_1ms_0/CS[7]_net_1 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_153 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m61  
        (.A(\s_acq_change_0_s_stripnum[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[1]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_2_i ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_62_i ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3_I_5  (
        .A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIIHJB2[0]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_3[1] ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[4]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[4] ));
    IOPAD_TRI \k1_pad/U0/U0  (.D(\k1_pad/U0/NET1 ), .E(
        \k1_pad/U0/NET2 ), .PAD(k1));
    NOR2B \scalestate_0/timecount_ret_38_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[3]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[3] ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[2]  (.D(
        \DUMP_0/dump_coder_0/para4_4[2]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[2]_net_1 ));
    DFN1 \CAL_0/cal_div_0/count[2]  (.D(\CAL_0/cal_div_0/count_5[2] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[2]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para3[11]  (.D(
        \DUMP_0/dump_coder_0/para4_4[11]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_4_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para3[11]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[23]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[23]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_299 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m49  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_46 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_49 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_50 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m136  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[3] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_137 ));
    DFN1 \timer_top_0/state_switch_0/dataout[8]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[8]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[8] ));
    DFN1 \state_1ms_0/timecount[16]  (.D(
        \state_1ms_0/timecount_RNO[16]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[16] ));
    NOR2B \s_acq_change_0/s_rst_RNO  (.A(\s_acq_change_0/N_68 ), .B(
        net_27), .Y(\s_acq_change_0/s_rst_RNO_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[6] ));
    MX2 \top_code_0/scan_rst_RNIQOT93  (.A(net_33), .B(\xa_c[0] ), .S(
        \top_code_0/N_258 ), .Y(\top_code_0/N_803 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m309  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_302 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_309 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[12] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_6_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_6_net ));
    IOTRI_OB_EB \Q4Q5_pad/U0/U1  (.D(Q4Q5_c), .E(VCC), .DOUT(
        \Q4Q5_pad/U0/NET1 ), .EOUT(\Q4Q5_pad/U0/NET2 ));
    DFN1E1 \plusestate_0/DUMPTIME[7]  (.D(\top_code_0_plusedata[7] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[7]_net_1 ));
    AND3 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2b_12_inst  
        (.A(\pd_pluse_top_0/count_6[3] ), .B(
        \pd_pluse_top_0/count_6[4] ), .C(\pd_pluse_top_0/count_1[5] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/incb_5_net )
        );
    XOR2 \PLUSE_0/bri_timer_0/count_RNO[5]  (.A(
        \PLUSE_0/bri_timer_0/count_c4 ), .B(\PLUSE_0/count_2[5] ), .Y(
        \PLUSE_0/bri_timer_0/count_n5 ));
    DFN1E1 \plusestate_0/PLUSETIME[9]  (.D(\top_code_0_plusedata[9] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[9]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNIDGCG[3]  (.A(
        \DUMP_0/dump_coder_0/para2[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_3[0] ));
    DFN1E1 \top_code_0/sd_sacq_data[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[3] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i22_mux ));
    DFN1E1 \scalestate_0/ACQ180_NUM[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[4]_net_1 ));
    XO1 \DUMP_0/dump_coder_0/para6_RNIOFI91[9]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_coder_0/para6[9]_net_1 ), .C(
        \DUMP_0/dump_coder_0/i_reg16_8[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_5[0] ));
    DFN1E1 \scanstate_0/acqtime[10]  (.D(\top_code_0_scandata[10] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[10]_net_1 ));
    OR3 \scalestate_0/timecount_ret_57_RNIS4I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[0] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[0] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[0] ), .Y(
        \scalestate_0_timecount[0] ));
    NOR2 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        );
    XOR2 \DUMP_0/dump_coder_0/para5_RNIIRLJ[4]  (.A(
        \DUMP_0/dump_coder_0/para5[4]_net_1 ), .B(\DUMP_0/count_1[4] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_0[0] ));
    DFN1E1 \scanstate_0/timecount_1[1]  (.D(
        \scanstate_0/timecount_5[1] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[1] ));
    XO1 \CAL_0/cal_div_0/count_RNI2KU71[5]  (.A(
        \CAL_0/cal_para_out[5] ), .B(\CAL_0/cal_div_0/count[5]_net_1 ), 
        .C(\CAL_0/cal_div_0/clear_n4_4 ), .Y(
        \CAL_0/cal_div_0/clear_n4_NE_0 ));
    XO1 \PLUSE_0/qq_coder_0/i_reg10_NE_0[0]  (.A(\PLUSE_0/count_9[4] ), 
        .B(\PLUSE_0/qq_para3[4] ), .C(\PLUSE_0/qq_para3[5] ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_NE_0[0]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[21]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[21]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_511 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/VXOR2_13_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_16_net ), 
        .B(\sd_acq_top_0/count[16] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[16] ));
    DFN1E1 \state_1ms_0/PLUSETIME[11]  (.D(
        \top_code_0_state_1ms_data[11] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[11]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[12]_net_1 ));
    AO1C \scalestate_0/necount_cmp_0/AO1C_0  (.A(
        \scalestate_0/necount[1]_net_1 ), .B(
        \scalestate_0/M_NUM[1]_net_1 ), .C(
        \scalestate_0/necount[0]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/AO1C_0_Y ));
    AO1 \state_1ms_0/timecount_RNO_2[13]  (.A(
        \state_1ms_0/M_DUMPTIME[13]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[13] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[13] ));
    OR2 \scalestate_0/CS_RNIPDHJ[8]  (.A(\scalestate_0/CS[8]_net_1 ), 
        .B(\scalestate_0/CS[9]_net_1 ), .Y(\scalestate_0/N_297 ));
    MX2C \DUMP_0/off_on_state_0/cs_RNO_0[1]  (.A(
        \DUMP_0/off_on_state_0/cs[1]_net_1 ), .B(\DUMP_0/i_1[1] ), .S(
        DUMP_0_dump_off), .Y(\DUMP_0/off_on_state_0/N_10 ));
    NOR2 \scalestate_0/timecount_ret_0_RNO  (.A(\scalestate_0/N_1206 ), 
        .B(\scalestate_0/un1_CS_20 ), .Y(
        \scalestate_0/timecount_cnst_m_0[6] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIPE8D[12]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[12]_net_1 )
        , .B(\pd_pluse_top_0/count[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_12[0] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_39_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m43_0 ));
    XO1 \DUMP_0/dump_coder_0/para5_RNIM9C71[9]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_coder_0/para5[9]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_5[0] ));
    DFN1 \DUMP_0/off_on_timer_1/count[0]  (.D(
        \DUMP_0/off_on_timer_1/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[0] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m221  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_222 ));
    DFN1E1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[2]  
        (.D(\top_code_0_s_periodnum[2] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[2]_net_1 )
        );
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m2_e  (.A(
        \top_code_0_s_addchoice[0] ), .B(\top_code_0_s_addchoice[1] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_311 ));
    DFN1E1 \top_code_0/scaleddsdiv[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[0] ));
    NOR2A \scalestate_0/CS_RNIJG2J[13]  (.A(\scalestate_0/N_1195 ), .B(
        \scalestate_0/CS[13]_net_1 ), .Y(\scalestate_0/N_1251_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[7]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[7] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[7]_net_1 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i2_mux ));
    NOR2 \top_code_0/s_acqnum_1_sqmuxa_0_a2_1  (.A(\top_code_0/N_150 ), 
        .B(\top_code_0/N_147 ), .Y(\top_code_0/s_acqnum_1_sqmuxa_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m177  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_176 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_177 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_178 ));
    DFN1E1 \scalestate_0/timecount_ret_41  (.D(
        \scalestate_0/timecount_20_iv_8[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[2] ));
    DFN1 \scalestate_0/dds_conf  (.D(
        \scalestate_0/dds_conf_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_dds_conf));
    MX2 \state_1ms_0/timecount_RNO_0[7]  (.A(
        \state_1ms_0/timecount_8[7] ), .B(\state_1ms_0_timecount[7] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_74 ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNI9FU2[4]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c2 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c4 ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[1]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs_i[0]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[1] ));
    MX2 \scalestate_0/strippluse_RNO_2[3]  (.A(
        \scalestate_0/STRIPNUM180_NUM[3]_net_1 ), .B(
        \scalestate_0/STRIPNUM90_NUM[3]_net_1 ), .S(
        \scalestate_0/N_1209_0 ), .Y(\scalestate_0/N_423 ));
    XNOR2 \scalestate_0/necount_cmp_0/XNOR2_8  (.A(
        \scalestate_0/necount[6]_net_1 ), .B(
        \scalestate_0/M_NUM[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/XNOR2_8_Y ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[0]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[0]_net_1 )
        );
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[4]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[8]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[7] ), 
        .Y(\DDS_0/dds_state_0/N_282 ));
    NOR3B \bridge_div_0/count_RNIJROM7[5]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[5]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIJROM7[5]_net_1 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[2]  (.D(
        \top_code_0_state_1ms_data[2] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[2]_net_1 ));
    NOR3B \scalestate_0/ACQ90_NUM_1_sqmuxa_0_a2  (.A(
        \scalestate_0/N_67 ), .B(\scalestate_0/N_62 ), .C(
        \top_code_0_scalechoice_0[0] ), .Y(
        \scalestate_0/ACQ90_NUM_1_sqmuxa ));
    DFN1 \scalestate_0/necount_LE_NE  (.D(
        \scalestate_0/necount_LE_NE_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        scalestate_0_ne_le));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_4  (.A(
        \scalestate_0/necount[10]_net_1 ), .B(
        \scalestate_0/NE_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_4_Y ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[10]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c8 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n10 ));
    AOI1B \DUMP_0/off_on_state_1/state_over_RNO_0  (.A(
        \DUMP_0/off_on_state_1/N_42_i ), .B(
        \DUMP_0/off_on_state_1_state_over ), .C(\DUMP_0/i_0[0] ), .Y(
        \DUMP_0/off_on_state_1/N_12_mux ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[17]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[18]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_500 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[4]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[5]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_318 ));
    XOR2 \DUMP_0/dump_coder_0/i_RNO_14[3]  (.A(
        \DUMP_0/dump_coder_0/para1[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_4_5[0] ));
    OA1C \top_code_0/state_1ms_load_RNO  (.A(\top_code_0/N_197 ), .B(
        top_code_0_state_1ms_load), .C(\top_code_0/N_314 ), .Y(
        \top_code_0/N_106 ));
    DFN1E1 \scalestate_0/timecount_ret_93  (.D(
        \scalestate_0/timecount_m3_e_2 ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_m3_e_2_reto ));
    DFN1 \scalestate_0/s_acqnum_1[4]  (.D(
        \scalestate_0/s_acqnum_1_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[4] ));
    OA1A \scalestate_0/necount_cmp_0/OA1A_0  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/M_NUM[9]_net_1 ), .C(
        \scalestate_0/M_NUM[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OA1A_0_Y ));
    MX2 \top_code_0/state_1ms_rst_n_0_0_RNIC5PK5  (.A(
        top_code_0_state_1ms_rst_n_0), .B(\top_code_0/un1_xa_2 ), .S(
        \top_code_0/N_320 ), .Y(\top_code_0/N_800 ));
    NOR3B \top_code_0/s_addchoice_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/s_addchoice_1_sqmuxa_0_a2_0_net_1 ), .C(
        \top_code_0/N_152 ), .Y(\top_code_0/s_addchoice_1_sqmuxa ));
    AO1C \state_1ms_0/CS_RNO_0[8]  (.A(\state_1ms_0/CS[7]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[8] ));
    NOR2B \top_code_0/relay_close_RNO[5]  (.A(\top_code_0/N_824 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[5]_net_1 ));
    DFN1 \top_code_0/relay_close[6]  (.D(
        \top_code_0/relay_close_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[6] ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[4] ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[10]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[10] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_1[10] ));
    AO1 \scalestate_0/timecount_ret_20_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[8]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[8] ), .Y(
        \scalestate_0/timecount_20_iv_4[8] ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[3]  (.A(
        \DDS_0/dds_state_0/para[3]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_489 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[3] ));
    AO1A \top_code_0/scale_start_ret_3_RNO  (.A(\top_code_0/N_174 ), 
        .B(\top_code_0/N_329 ), .C(\top_code_0/N_162 ), .Y(
        \top_code_0/N_110 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[11]_net_1 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_13  (.A(\xd_in[1] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[1] ));
    AO1 \scalestate_0/timecount_ret_47_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[16]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[16] ), .Y(
        \scalestate_0/timecount_20_0_iv_2[16] ));
    OR3 \top_code_0/s_load_3_i_o2  (.A(\xa_c[6] ), .B(
        \top_code_0/N_137 ), .C(\top_code_0/N_140 ), .Y(
        \top_code_0/N_152 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[6]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[6] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[6] ));
    IOPAD_TRI \pulse_start_pad/U0/U0  (.D(\pulse_start_pad/U0/NET1 ), 
        .E(\pulse_start_pad/U0/NET2 ), .PAD(pulse_start));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[0]  (.A(
        \scalestate_0/ACQ180_NUM[0]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[0]_net_1 ), .S(\scalestate_0/N_1209_0 )
        , .Y(\scalestate_0/N_448 ));
    DFN1 \s_acq_change_0/s_acqnum[1]  (.D(
        \s_acq_change_0/s_acqnum_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[1] ));
    OR3 \DUMP_0/dump_coder_0/para6_RNIKOPR2[6]  (.A(
        \DUMP_0/dump_coder_0/i_reg16_7[0] ), .B(
        \DUMP_0/dump_coder_0/i_reg16_11[0] ), .C(
        \DUMP_0/dump_coder_0/i_reg16_NE_1[0] ), .Y(
        \DUMP_0/dump_coder_0/i_reg16_NE_6[0] ));
    IOPAD_IN \xwe_pad/U0/U0  (.PAD(xwe), .Y(\xwe_pad/U0/NET1 ));
    DFN1 \scalestate_0/necount[8]  (.D(
        \scalestate_0/necount_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0/necount[8]_net_1 ));
    NOR2A \pd_pluse_top_0/pd_pluse_coder_0/i_RNO[2]  (.A(net_27), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_1[2] ));
    DFN1 \DUMP_0/dump_state_0/cs[4]  (.D(
        \DUMP_0/dump_state_0/cs_RNO_0[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[4]_net_1 ));
    IOTRI_OR_EB \ddsreset_pad/U0/U1  (.D(
        \DDS_0/dds_state_0/reset_RNO_net_1 ), .E(VCC), .OCLK(GLA_net_1)
        , .DOUT(\ddsreset_pad/U0/NET1 ), .EOUT(\ddsreset_pad/U0/NET2 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m305  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[12] ), .C(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_306 ));
    OR2A \PLUSE_0/qq_state_0/cs_RNO_0[1]  (.A(
        \PLUSE_0/qq_state_0/cs[1]_net_1 ), .B(\PLUSE_0/i_9[1] ), .Y(
        \PLUSE_0/qq_state_0/N_82 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m45_0 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_1_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_6_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_1_net ));
    NOR2B \state_1ms_0/timecount_RNO_5[13]  (.A(
        \state_1ms_0/PLUSECYCLE[13]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[13] ));
    DFN1E1 \scalestate_0/M_NUM[10]  (.D(\top_code_0_scaledatain[10] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[10]_net_1 ));
    NOR2B \DDS_0/dds_state_0/reset_RNO  (.A(
        \DDS_0/dds_state_0/cs[1]_net_1 ), .B(\DDS_0/dds_state_0/N_223 )
        , .Y(\DDS_0/dds_state_0/reset_RNO_net_1 ));
    OA1 \ClockManagement_0/long_timer_0/timeup_RNO  (.A(sigtimeup_c), 
        .B(\ClockManagement_0/long_timer_0/timeup_0_sqmuxa ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_RNO_net_1 ));
    DFN1 \top_code_0/relay_on[8]  (.D(
        \top_code_0/relay_on_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[8] ));
    NOR2A \scalestate_0/ACQTIME_1_sqmuxa_0_a2_0  (.A(
        \top_code_0_scalechoice_0[3] ), .B(
        \top_code_0_scalechoice_0[2] ), .Y(\scalestate_0/N_65 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m44_0 ));
    XO1 \scalestate_0/fst_lst_pulse_RNO_2  (.A(
        \scalestate_0/necount[4]_net_1 ), .B(
        \scalestate_0/NE_NUM[4]_net_1 ), .C(
        \scalestate_0/fst_lst_pulse8_10 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_4 ));
    AND3 \bridge_div_0/count_5_I_10  (.A(
        \bridge_div_0/count_RNIEMOM7[0]_net_1 ), .B(
        \bridge_div_0/count_RNIFNOM7[1]_net_1 ), .C(
        \bridge_div_0/count_RNIGOOM7[2]_net_1 ), .Y(
        \bridge_div_0/DWACT_FINC_E[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[14]  (.A(
        \state_1ms_0_timecount[14] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_262 ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[5] ));
    NOR2A \scalestate_0/timecount_ret_56_RNO_3  (.A(
        \scalestate_0/CUTTIME90[19]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[19] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_143  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_76_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_51_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_143_Y ));
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_RNO  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_net_1 ), 
        .B(n_acq_change_0_n_rst_n), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_RNO_net_1 )
        );
    AO1A \scalestate_0/timecount_ret_10_RNIO241  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .B(
        \scalestate_0/timecount_cnst_m_0_reto[7] ), .C(
        \scalestate_0/timecount_20_iv_10_reto[7] ), .Y(
        \scalestate_0_timecount[7] ));
    NOR2B \scalestate_0/necount_RNO[5]  (.A(\scalestate_0/N_735 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[5]_net_1 ));
    DFN1 \topctrlchange_0/rt_sw  (.D(\topctrlchange_0/rt_sw_RNO_4 ), 
        .CLK(GLA_net_1), .Q(rt_sw_net_0));
    NOR2B \state_1ms_0/timecount_RNO[17]  (.A(\state_1ms_0/N_84 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[17]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME90[6]  (.D(\top_code_0_scaledatain[6] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1685 ), .Q(
        \scalestate_0/CUTTIME90[6]_net_1 ));
    OA1C \scalestate_0/necount_cmp_1/OA1C_0  (.A(
        \scalestate_0/necount[9]_net_1 ), .B(
        \scalestate_0/NE_NUM[9]_net_1 ), .C(
        \scalestate_0/necount[10]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/OA1C_0_Y ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[23]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[23]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_300 ));
    DFN1E1 \state_1ms_0/PLUSETIME[6]  (.D(
        \top_code_0_state_1ms_data[6] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[6]_net_1 ));
    MX2 \scan_scale_sw_0/s_start_RNO_1  (.A(scanstate_0_s_acq), .B(
        sd_acq_en_c), .S(\top_code_0_change_0[0] ), .Y(
        \scan_scale_sw_0/s_start_5 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m156  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_155 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_156 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_157 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_64  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_64_Y ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNIMEEH[10]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[10]_net_1 )
        , .B(\pd_pluse_top_0/count_0[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_10[0] ));
    MX2 \noisestate_0/timecount_1_RNO_0[5]  (.A(
        \noisestate_0/acqtime[5]_net_1 ), .B(
        \noisestate_0/dectime[5]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_62 ));
    OR3 \DUMP_0/dump_coder_0/para4_RNIOLAA2[2]  (.A(
        \DUMP_0/dump_coder_0/un1_count_1_3[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_4[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_1_NE_3[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_7[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[1]  (.D(
        \DUMP_0/dump_coder_0/para2_4[1]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[1]_net_1 ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_0  (.A(
        \scalestate_0/necount_cmp_0/NOR3A_0_Y ), .B(
        \scalestate_0/necount_cmp_0/OR2A_5_Y ), .C(
        \scalestate_0/necount_cmp_0/NAND3A_2_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_0_Y ));
    DFN1 \top_code_0/scale_start_ret  (.D(top_code_0_scale_start), 
        .CLK(GLA_net_1), .Q(\top_code_0/top_code_0_scale_start_reto ));
    DFN1E1 \top_code_0/n_divnum[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[8] ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[11]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[11] ), .CLK(ddsclkout_c)
        , .Q(\sd_acq_top_0/sd_sacq_state_0/cs[11]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[2]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[2]_net_1 ));
    NOR3A \top_code_0/un1_xa_8_16_i_i_o3_i_a2_4  (.A(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_1_net_1 ), .B(\xa_c[11] ), 
        .C(\xa_c[12] ), .Y(
        \top_code_0/un1_xa_8_16_i_i_o3_i_a2_4_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[1]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_14_i ), .CLK(
        GLA_net_1), .E(top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[1]_net_1 ));
    AO1A \scalestate_0/timecount_ret_34_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[9]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[9] ), .Y(
        \scalestate_0/timecount_20_iv_1[9] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[13]  (.D(
        \top_code_0_dds_configdata[12] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[13]_net_1 ));
    DFN1E1 \scalestate_0/timecount_ret_61  (.D(
        \scalestate_0/timecount_20_iv_6[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[12] ));
    XA1 \PLUSE_0/qq_timer_0/count_RNO[3]  (.A(
        \PLUSE_0/qq_timer_0/count_c2 ), .B(\PLUSE_0/count_9[3] ), .C(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_0/count_n3 ));
    OA1C \PLUSE_0/qq_state_1/cs_RNO_0[2]  (.A(Q4Q5_c), .B(
        \PLUSE_0/i_2[2] ), .C(\PLUSE_0/qq_state_1/cs[1]_net_1 ), .Y(
        \PLUSE_0/qq_state_1/N_89 ));
    XA1 \PLUSE_0/qq_timer_1/count_RNO[4]  (.A(
        \PLUSE_0/qq_timer_1/count_9_0 ), .B(\PLUSE_0/count_7[4] ), .C(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_1/count_n4 ));
    DFN1E1 \top_code_0/n_divnum[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[2] ));
    RAM512X18 #( .MEMORYFILE("RAM_R4C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R4C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_4_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_4_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_0_net ));
    DFN1 \noisestate_0/CS[1]  (.D(\noisestate_0/CS_RNO[1]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[1]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_59  (.A(
        \timer_top_0/timer_0/N_3 ), .B(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .Y(
        \timer_top_0/timer_0/I_59 ));
    XA1A \timer_top_0/timer_0/Timer_Cmp_0/AND2_1  (.A(
        \timer_top_0/dataout[21] ), .B(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_9_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_1_Y ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[5]  (.D(
        \top_code_0_pd_pluse_data[5] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[5]_net_1 ));
    NOR3C \ClockManagement_0/long_timer_0/count_RNIHHP03[3]  (.A(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_2 ), .B(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_1 ), .C(
        \ClockManagement_0/long_timer_0/count_c2 ), .Y(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_7 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIF1LR[3]  (.A(
        \ClockManagement_0/long_timer_0/count[3]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[4]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_1 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_1_12_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_5_net ), 
        .C(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ));
    OR3 \DDS_0/dds_state_0/para_RNO[7]  (.A(\DDS_0/dds_state_0/N_273 ), 
        .B(\DDS_0/dds_state_0/N_272 ), .C(
        \DDS_0/dds_state_0/para_9_i_i_1[7] ), .Y(
        \DDS_0/dds_state_0/N_8 ));
    IOIN_IB \ADC_pad[5]/U0/U1  (.YIN(\ADC_pad[5]/U0/NET1 ), .Y(
        \ADC_c[5] ));
    RAM512X18 #( .MEMORYFILE("RAM_R12C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R12C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_12_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_12_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_0_net )
        );
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI4B09[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_22[0] ));
    MX2 \plusestate_0/timecount_1_RNO_0[15]  (.A(
        \plusestate_0/DUMPTIME[15]_net_1 ), .B(
        \plusestate_0/PLUSETIME[15]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_86 ));
    DFN1 \noisestate_0/dumpon_ctr  (.D(
        \noisestate_0/dumpon_ctr_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        noisestate_0_dumpon_ctr));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m174  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_159 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_174 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[2] ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_15[10]  (.A(
        \sd_acq_top_0/count_3[7] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[7]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_6[10] ));
    NOR3C \top_code_0/pluse_str_RNO_1  (.A(\top_code_0/N_339 ), .B(
        \top_code_0/N_336 ), .C(\top_code_0/un1_xa_49_0_a2_1 ), .Y(
        \top_code_0/un1_xa_49 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_4  (.A(
        \timer_top_0/dataout[4] ), .B(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_10_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_4_Y ));
    DFN1 \s_acq_change_0/s_acqnum[13]  (.D(
        \s_acq_change_0/s_acqnum_RNO[13]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[13] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIDS6T[18]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[18]_net_1 ), .B(
        \sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_18[0] ));
    AX1C \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/POR2_9_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net )
        , .C(\pd_pluse_top_0/count[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[12] ));
    DFN1E1 \scalestate_0/timecount_ret_53  (.D(
        \scalestate_0/timecount_20_0_iv_4[18] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_4_reto[18] ));
    XOR2 \scalestate_0/M_pulse_RNO_14  (.A(
        \scalestate_0/M_NUM[9]_net_1 ), .B(
        \scalestate_0/necount[9]_net_1 ), .Y(\scalestate_0/M_pulse8_9 )
        );
    MX2A \plusestate_0/sw_acq1_RNO_0  (.A(\plusestate_0/N_302 ), .B(
        plusestate_0_sw_acq1), .S(\plusestate_0/N_298 ), .Y(
        \plusestate_0/N_120 ));
    DFN1E1 \state_1ms_0/CUTTIME[18]  (.D(
        \top_code_0_state_1ms_data[2] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_380 ), .Q(\state_1ms_0/CUTTIME[18]_net_1 ));
    XOR2 \PLUSE_0/qq_coder_0/un1_qq_para2_0[0]  (.A(
        \PLUSE_0/qq_para2[0] ), .B(\PLUSE_0/count_9[0] ), .Y(
        \PLUSE_0/qq_coder_0/un1_qq_para2_0[0]_net_1 ));
    DFN1 \DUMP_OFF_1/off_on_state_0/state_over  (.D(
        \DUMP_OFF_1/off_on_state_0/N_9 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/off_on_state_0_state_over ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m100  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_99 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_100 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_101 ));
    OR3 \scalestate_0/timecount_ret_1_RNO  (.A(
        \scalestate_0/timecount_20_iv_3[5] ), .B(
        \scalestate_0/timecount_20_iv_2[5] ), .C(
        \scalestate_0/timecount_20_iv_6[5] ), .Y(
        \scalestate_0/timecount_20_iv_9[5] ));
    XOR2 \PLUSE_0/qq_coder_1/i_RNO_3[1]  (.A(\PLUSE_0/qq_para1[1] ), 
        .B(\PLUSE_0/count_7[1] ), .Y(
        \PLUSE_0/qq_coder_1/un1_count_1[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[7]  (.D(
        \DUMP_0/dump_coder_0/para4_4[7]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[7]_net_1 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[1]_net_1 ));
    NOR2A \scalestate_0/timecount_ret_67_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[14]_net_1 ), .B(\scalestate_0/N_1089 )
        , .Y(\scalestate_0/S_DUMPTIME_m[14] ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[0]  (.D(
        \top_code_0_cal_data[0] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[0] ));
    DFN1E1 \noisestate_0/acqtime[5]  (.D(\top_code_0_noisedata[5] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[5]_net_1 ));
    NOR2B \state_1ms_0/bri_cycle_RNO  (.A(\state_1ms_0/N_156 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/bri_cycle_RNO_0_net_1 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m36  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[12]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[13]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i22_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_37_i ));
    NOR3B \bridge_div_0/count_RNIGOOM7[2]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[2]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIGOOM7[2]_net_1 ));
    AO1A \scalestate_0/timecount_20_iv_5_RNO[5]  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[5]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[5] ), .Y(
        \scalestate_0/timecount_20_iv_0[5] ));
    XO1 \scalestate_0/fst_lst_pulse_RNO_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/NE_NUM[8]_net_1 ), .C(
        \scalestate_0/fst_lst_pulse8_7 ), .Y(
        \scalestate_0/fst_lst_pulse8_NE_3 ));
    DFN1 \PLUSE_0/qq_timer_0/count[2]  (.D(
        \PLUSE_0/qq_timer_0/count_n2 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_9[2] ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[8]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO_1[8] ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[8]_net_1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[1]  (.A(
        \s_acq_change_0/s_stripnum_5[1] ), .B(
        \s_acq_change_0_s_stripnum[1] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_57 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m290  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_291 ));
    DFN1E1 \top_code_0/sigtimedata[10]  (.D(\GPMI_0_dataout[10] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[10] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m37  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[0] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_38 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_135  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_128_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_47_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_135_Y ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_1_0 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I0_un1_CO1 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0 )
        );
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m41_3 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_116  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_98_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_27_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_116_Y ));
    OR3 \scalestate_0/timecount_ret_35_RNO_2  (.A(
        \scalestate_0/PLUSETIME180_m[9] ), .B(
        \scalestate_0/ACQTIME_m[9] ), .C(
        \scalestate_0/OPENTIME_TEL_m[9] ), .Y(
        \scalestate_0/timecount_20_iv_5[9] ));
    NOR3B \scalestate_0/M_NUM_1_sqmuxa_0_a2_1  (.A(
        top_code_0_scaleload), .B(\top_code_0_scalechoice_0[4] ), .C(
        \top_code_0_scalechoice_0[1] ), .Y(\scalestate_0/N_64 ));
    OR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_8  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[4]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_9 ));
    AX1C \ClockManagement_0/clk_10k_0/un1_count_1_I_37  (.A(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \ClockManagement_0/clk_10k_0/count[2]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/count[3]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/I_37_0 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_RNO_net_1 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk_net_1 ));
    NOR2B \top_code_0/noisedata_1_sqmuxa_0_a2_0_0  (.A(
        \top_code_0/N_333 ), .B(net_27), .Y(
        \top_code_0/noisedata_1_sqmuxa_0_a2_0_net_1 ));
    MX2 \plusestate_0/timecount_1_RNO_0[0]  (.A(
        \plusestate_0/DUMPTIME[0]_net_1 ), .B(
        \plusestate_0/PLUSETIME[0]_net_1 ), .S(\plusestate_0/N_213 ), 
        .Y(\plusestate_0/N_71 ));
    AND2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_15  
        (.A(\s_acq_change_0_s_stripnum[3] ), .B(
        \s_acq_change_0_s_stripnum[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[1] )
        );
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[2]  (.D(
        \top_code_0_pd_pluse_data[2] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[2]_net_1 ));
    IOIN_IB \xa_pad[11]/U0/U1  (.YIN(\xa_pad[11]/U0/NET1 ), .Y(
        \xa_c[11] ));
    NOR3B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_RNO[2]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_7_1 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[2] ));
    DFN1 \DUMP_OFF_0/off_on_coder_0/i[1]  (.D(
        \DUMP_OFF_0/off_on_coder_0/i_RNO_3[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/i_3[1] ));
    DFN1 \DDS_0/dds_timer_0/count[4]  (.D(\DDS_0/dds_timer_0/count_n4 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[4] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[2]  (.D(
        \top_code_0_state_1ms_data[2] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[2]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[17]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m42_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[17] ));
    OR2A \scanstate_0/sw_acq2_RNO  (.A(net_33), .B(\scanstate_0/N_109 )
        , .Y(\scanstate_0/sw_acq2_RNO_2 ));
    AO1C \state_1ms_0/CS_RNO_0[9]  (.A(\state_1ms_0/CS[8]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[9] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m193  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_194 ));
    NOR3 \top_code_0/n_load_RNO_1  (.A(\top_code_0/N_154 ), .B(
        \top_code_0/N_152 ), .C(\top_code_0/N_159 ), .Y(
        \top_code_0/N_280 ));
    XA1 \DDS_0/dds_timer_0/count_RNO[2]  (.A(
        \DDS_0/dds_timer_0/count_c1 ), .B(\DDS_0/count[2] ), .C(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DDS_0/dds_timer_0/count_n2 ));
    IOPAD_IN \zcs2_pad/U0/U0  (.PAD(zcs2), .Y(\zcs2_pad/U0/NET1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[3]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c2 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[3]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n3 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI85JS[2]  (.A(
        \sd_acq_top_0/count_10[2] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[2]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_6[0] ));
    NOR2A \scalestate_0/strippluse_RNO_1[8]  (.A(\scalestate_0/N_428 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[8] ));
    DFN1E1 \top_code_0/state_1ms_data[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[13] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[4] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_64_i ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa_0_a2  (
        .A(\top_code_0_sd_sacq_choice[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_3_i_a2_1 ), 
        .Y(\sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ));
    XA1A \PLUSE_0/qq_coder_1/i_RNO_2[1]  (.A(\PLUSE_0/count_7[0] ), .B(
        \PLUSE_0/qq_para1[0] ), .C(\PLUSE_0/qq_coder_1/i_0_0[1] ), .Y(
        \PLUSE_0/qq_coder_1/i_0_2[1] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m47_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_12  (.A(
        \scalestate_0/NE_NUM[0]_net_1 ), .B(
        \scalestate_0/necount[0]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_0 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m13  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[1] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_14_0 ));
    DFN1C0 \syn_md_module_1/syn_md_edge_detect_0/sig_r0  (.D(
        syn_md_tmp_c), .CLK(GLA_net_1), .CLR(top_code_0_scale_rst_0), 
        .Q(\syn_md_module_1/syn_md_edge_detect_0/sig_r0_net_1 ));
    AO1 \scalestate_0/timecount_ret_53_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[18]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[18] ), .Y(
        \scalestate_0/timecount_20_0_iv_2[18] ));
    NOR2B \scalestate_0/strippluse_RNO[11]  (.A(\scalestate_0/N_570 ), 
        .B(top_code_0_scale_rst_3), .Y(
        \scalestate_0/strippluse_RNO[11]_net_1 ));
    NOR2B \DUMP_0/off_on_timer_1/count_RNIJQ3N[1]  (.A(
        \DUMP_0/count_0[0] ), .B(\DUMP_0/count_0[1] ), .Y(
        \DUMP_0/off_on_timer_1/count_c1 ));
    AO1A \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNO  (
        .A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_i ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNO_net_1 )
        );
    NOR2B \top_code_0/relay_close_RNO[1]  (.A(\top_code_0/N_820 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[1]_net_1 ));
    AO1 \scalestate_0/timecount_RNO_0[20]  (.A(
        \scalestate_0/CUTTIME180_TEL[20]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[20] )
        , .Y(\scalestate_0/timecount_20_0_iv_0[20] ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/TND2_15_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_16_net ), 
        .B(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_17_net )
        , .C(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_22_net ), 
        .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_15_net ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[5]_net_1 ));
    OR3 \DUMP_0/dump_coder_0/para3_RNI8HB52[11]  (.A(
        \DUMP_0/dump_coder_0/un1_count_2_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_2_11[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE_1[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_6[0] ));
    XOR2 \bridge_div_0/dataall_RNI4SNO[0]  (.A(
        \bridge_div_0/dataall[0]_net_1 ), .B(
        \bridge_div_0/count[0]_net_1 ), .Y(
        \bridge_div_0/un1_count_0[0] ));
    DFN1E1 \top_code_0/dds_configdata[8]  (.D(\GPMI_0_dataout[8] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[8] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m147  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_148 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[17]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[17]_net_1 ));
    DFN1 \timer_top_0/timer_0/timedata[20]  (.D(
        \timer_top_0/timer_0/timedata_4[20] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[20]_net_1 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[24]  (.A(
        \top_code_0_dds_configdata[7] ), .B(\DDS_0/dds_state_0/N_569 ), 
        .C(\DDS_0/dds_state_0/N_303 ), .Y(
        \DDS_0/dds_state_0/para_9_i_1[24] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[9]_net_1 ));
    NOR2A \scalestate_0/CS_RNO[13]  (.A(top_code_0_scale_rst_5), .B(
        \scalestate_0/N_1237 ), .Y(\scalestate_0/CS_RNO[13]_net_1 ));
    OR2 \scalestate_0/timecount_ret_17_RNI61C  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_1_reto ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_9_reto ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ));
    NOR3 \top_code_0/dump_sustain_RNO_1  (.A(\top_code_0/N_144 ), .B(
        \top_code_0/N_167 ), .C(\top_code_0/N_161 ), .Y(
        \top_code_0/N_262 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[16]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[16] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[16] ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[3]  (.D(
        \top_code_0_cal_data[3] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[3] ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_2  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_7_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_6_Y ), .C(
        \timer_top_0/dataout[15] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_2_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[1] ));
    AO1B \sd_acq_top_0/sd_sacq_state_0/stateover_RNO  (.A(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_245 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/stateover_RNO_2 ));
    DFN1 \PLUSE_0/qq_coder_1/i[2]  (.D(\PLUSE_0/qq_coder_1/i_RNO_3[2] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_2[2] ));
    NOR3C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[11]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/i_1[3] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs[10]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[11]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_41_RNO_3  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[2]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[2] ));
    DFN1 \state_1ms_0/rt_sw  (.D(\state_1ms_0/rt_sw_RNO_3 ), .CLK(
        GLA_net_1), .Q(state_1ms_0_rt_sw));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m135  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[19] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_136 ));
    NOR3B \top_code_0/state_1ms_data_1_sqmuxa_0_a2  (.A(net_27), .B(
        \top_code_0/state_1ms_data_1_sqmuxa_0_a2_1_net_1 ), .C(
        \top_code_0/N_152 ), .Y(\top_code_0/state_1ms_data_1_sqmuxa ));
    OR2A \scalestate_0/s_acq180_RNO_1  (.A(timer_top_0_clk_en_scale), 
        .B(\scalestate_0/un1_CS6_0 ), .Y(\scalestate_0/un1_CS6 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i8_mux ));
    AX1C \ClockManagement_0/clk_div500_0/un1_count_1_I_38  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] ), 
        .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_2[0] )
        , .C(\ClockManagement_0/clk_div500_0/count[8]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/I_38 ));
    IOPAD_BI \xd_pad[1]/U0/U0  (.D(\xd_pad[1]/U0/NET1 ), .E(
        \xd_pad[1]/U0/NET2 ), .Y(\xd_pad[1]/U0/NET3 ), .PAD(xd[1]));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[6]_net_1 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[8]  (.A(
        \timer_top_0/state_switch_0/N_247 ), .B(
        \timer_top_0/state_switch_0/N_249 ), .C(
        \timer_top_0/state_switch_0/N_248 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[8] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_5  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_164_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_79_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_5_Y ));
    OR2 \top_code_0/un1_state_1ms_rst_n117_4_i_o2_0  (.A(
        \top_code_0/N_139 ), .B(\xa_c[7] ), .Y(\top_code_0/N_171 ));
    OA1B \top_code_0/pluse_noise_ctrl_RNO_0  (.A(\xa_c[1] ), .B(
        \top_code_0/N_176 ), .C(top_code_0_pluse_noise_ctrl), .Y(
        \top_code_0/N_293 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[18]  (.A(
        \scalestate_0_timecount[18] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_270 ));
    NOR3 \scalestate_0/necount_cmp_1/NOR3_0  (.A(
        \scalestate_0/necount_cmp_1/OA1A_0_Y ), .B(
        \scalestate_0/necount_cmp_1/AND2A_0_Y ), .C(
        \scalestate_0/necount_cmp_1/OA1C_0_Y ), .Y(
        \scalestate_0/necount_cmp_1/NOR3_0_Y ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[0] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_2_i ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNIGPLJ[3]  (.A(
        \DUMP_0/dump_coder_0/para5[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_0[0] ));
    DFN1E1 \top_code_0/scaleddsdiv[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaleddsdiv_1_sqmuxa ), .Q(
        \top_code_0_scaleddsdiv[2] ));
    DFN1E1 \top_code_0/sigtimedata[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[4] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_0_RNO  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[0]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[0]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_0_i_i )
        );
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_15  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m38 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[0] )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i14_mux ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[1]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(\top_code_0_dds_configdata[0] ), 
        .Y(\DDS_0/dds_state_0/N_278 ));
    IOIN_IB \ADC_pad[6]/U0/U1  (.YIN(\ADC_pad[6]/U0/NET1 ), .Y(
        \ADC_c[6] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_50  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_145_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_97_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_50_Y ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[9]_net_1 ));
    DFN1E1 \top_code_0/scandata[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[8] ));
    DFN1E1 \top_code_0/sd_sacq_data[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[14] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m180  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_179 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_180 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_181 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[7]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[7] ));
    NOR2A \s_acq_change_0/s_acqnum_RNO_1[13]  (.A(
        \top_code_0_s_acqnum_2[13] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[13] ));
    MX2 \scanstate_0/timecount_1_RNO_0[5]  (.A(
        \scanstate_0/acqtime[5]_net_1 ), .B(
        \scanstate_0/dectime[5]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_63 ));
    AO1B \pd_pluse_top_0/pd_pluse_state_0/stateover_RNO  (.A(
        \pd_pluse_top_0/pd_pluse_state_0_stateover ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_195 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/stateover_RNO_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[6]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[6] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m266  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_267 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_3_inst  (.A(
        \sd_acq_top_0/count_10[0] ), .B(\sd_acq_top_0/count_10[1] ), 
        .C(\sd_acq_top_0/count_10[2] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ));
    DFN1E1 \scalestate_0/timecount_ret_25  (.D(
        \scalestate_0/timecount_20_iv_3[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_3_reto[11] ));
    IOPAD_IN \ADC_pad[11]/U0/U0  (.PAD(ADC[11]), .Y(
        \ADC_pad[11]/U0/NET1 ));
    NOR2B \state_1ms_0/timecount_RNO_5[3]  (.A(
        \state_1ms_0/PLUSETIME[3]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m70_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[0] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[1]  (.D(
        \top_code_0_n_divnum_0[1] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[1]_net_1 ));
    OR2 \scalestate_0/timecount_ret_10_RNO_0  (.A(
        \scalestate_0/CS[13]_net_1 ), .B(
        \scalestate_0/timecount_11_sqmuxa ), .Y(
        \scalestate_0/N_508_i_0_0 ));
    DFN1E1 \scanstate_0/acqtime[12]  (.D(\top_code_0_scandata[12] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[12]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[12]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[12]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_332 ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[11]  (.A(
        \top_code_0_dumpdata_0[11] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[11] ));
    NOR2A \DDS_0/dds_state_0/para_9_i_0_a2_4_0[22]  (.A(\DDS_0/i[0] ), 
        .B(top_code_0_dds_load), .Y(\DDS_0/dds_state_0/N_534_0 ));
    MX2 \scanstate_0/timecount_1_RNO[2]  (.A(\scanstate_0/N_60 ), .B(
        \scanstate_0/timecount_cnst[2] ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[2] ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[3]  (.D(
        \ClockManagement_0/long_timer_0/count_n3 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[3]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m51  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[16] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_52 ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_10  (.A(
        \timer_top_0/dataout[18] ), .B(
        \timer_top_0/timer_0/timedata[18]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_6_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_10_Y ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m70  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m70_3 ));
    XA1 \DUMP_OFF_1/off_on_timer_0/count_RNO[3]  (.A(
        \DUMP_OFF_1/off_on_timer_0/count_c2 ), .B(
        \DUMP_OFF_1/count_4[3] ), .C(
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_n3 ));
    OR2 \top_code_0/scaleload_3_i_o2  (.A(\top_code_0/N_148 ), .B(
        \top_code_0/N_150 ), .Y(\top_code_0/N_174 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_62_i ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[13]  (.A(
        \scanstate_0_timecount[13] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_191 ));
    DFN1E1 \top_code_0/scaledatain_0[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain_0[3] ));
    AO1A \scalestate_0/timecount_ret_20_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[8]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[8] ), .Y(
        \scalestate_0/timecount_20_iv_0[8] ));
    DFN1C0 \PLUSE_0/bri_coder_0/i[1]/U1  (.D(
        \PLUSE_0/bri_coder_0/i[1]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/i_8[1] ));
    DFN1 \scalestate_0/strippluse[3]  (.D(
        \scalestate_0/strippluse_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[3] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_1  
        (.A(\s_acq_change_0_s_stripnum[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I10_un1_CO1 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_12 )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_148  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_64_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_114_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_148_Y ));
    DFN1E1 \scanstate_0/acqtime[4]  (.D(\top_code_0_scandata[4] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[4]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[11]_net_1 ));
    DFN1 \timer_top_0/timer_0/timedata[21]  (.D(
        \timer_top_0/timer_0/timedata_4[21] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[21]_net_1 ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[6]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[6] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[5]  (.A(
        \plusestate_0_timecount[5] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_219 ));
    MX2 \scalestate_0/necount_RNO_0[7]  (.A(\scalestate_0/necount1[7] )
        , .B(\scalestate_0/necount[7]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_737 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m122  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_121 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_122 ), .S(
        \top_code_0_s_addchoice_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_123 ));
    NOR2B \DDS_0/dds_state_0/cs_RNO[6]  (.A(
        \DDS_0/dds_state_0/cs[5]_net_1 ), .B(\DDS_0/dds_state_0/N_223 )
        , .Y(\DDS_0/dds_state_0/cs_RNO[6]_net_1 ));
    AX1C \ClockManagement_0/clk_div500_0/un1_count_1_I_32  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_2[0] ), 
        .B(\ClockManagement_0/clk_div500_0/count[4]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count[5]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/I_32 ));
    NOR3C \ClockManagement_0/clk_10k_0/un1_count_1_I_43  (.A(
        \ClockManagement_0/clk_10k_0/count[2]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[3]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_1[0] ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_2[0] ));
    IOPAD_TRI \relay_close_pad[3]/U0/U0  (.D(
        \relay_close_pad[3]/U0/NET1 ), .E(\relay_close_pad[3]/U0/NET2 )
        , .PAD(relay_close[3]));
    IOIN_IB \xa_pad[12]/U0/U1  (.YIN(\xa_pad[12]/U0/NET1 ), .Y(
        \xa_c[12] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataeight[7]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataeight_1_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[7] ));
    IOPAD_TRI \relay_close_pad[4]/U0/U0  (.D(
        \relay_close_pad[4]/U0/NET1 ), .E(\relay_close_pad[4]/U0/NET2 )
        , .PAD(relay_close[4]));
    DFN1E1 \top_code_0/scandata[13]  (.D(\GPMI_0_dataout[13] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[13] ));
    NOR2 \state_1ms_0/dump_start_RNO_2  (.A(\state_1ms_0/CS[2]_net_1 ), 
        .B(\state_1ms_0/CS[7]_net_1 ), .Y(
        \state_1ms_0/un1_CS_9_0_a4_0 ));
    NOR3A \DUMP_0/dump_coder_0/i_RNO_4[3]  (.A(
        \DUMP_0/dump_coder_0/i_0_0_a2_5[3] ), .B(
        \DUMP_0/dump_coder_0/un1_count_4_8[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_4_9[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_8[3] ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/ADD_20x20_slow_I19_Y_2 )
        );
    DFN1E1 \scalestate_0/OPENTIME[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[10]_net_1 ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7_RNI8HLJ  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_8_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7_net_1 )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIDM3A[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_9[0] ));
    NOR2B \scalestate_0/timecount_ret_5_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[2]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[2] ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[3]  (.A(\scalestate_0/N_550 ), 
        .B(top_code_0_scale_rst_5), .Y(
        \scalestate_0/s_acqnum_1_RNO[3]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_37_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[3]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[3] ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[9]  (.A(
        \s_acq_change_0/s_stripnum_5[9] ), .B(
        \s_acq_change_0_s_stripnum[9] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_65 ));
    DFN1E1 \top_code_0/n_acqnum[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[7] ));
    NOR2B \DUMP_0/off_on_coder_0/i_RNO[0]  (.A(
        \DUMP_0/dump_state_0_on_start ), .B(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_coder_0/i_RNO_2[0] ));
    OR3 \timer_top_0/state_switch_0/state_start_RNO_0  (.A(
        \timer_top_0/state_switch_0/N_289 ), .B(
        \timer_top_0/state_switch_0/N_297 ), .C(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/state_start5_0_0_1 ));
    XAI1 \scalestate_0/necount_RNO[0]  (.A(\scalestate_0/N_1179 ), .B(
        \scalestate_0/necount[0]_net_1 ), .C(top_code_0_scale_rst_4), 
        .Y(\scalestate_0/necount_RNO[0]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m168  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_167 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_168 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_169 ));
    OR2A \scalestate_0/CS_RNI2T6K1[21]  (.A(\scalestate_0/N_1209 ), .B(
        \scalestate_0/N_1201 ), .Y(\scalestate_0/N_1153_1 ));
    DFN1E1 \top_code_0/noisedata[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[0] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[10]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c9 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[10] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n10 ));
    AX1C \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_2_1_inst  (
        .A(\sd_acq_top_0/count_10[0] ), .B(\sd_acq_top_0/count_10[1] ), 
        .C(\sd_acq_top_0/count_10[2] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[2] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i16_mux ));
    NOR2A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[8]  (.A(net_27), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[8] ));
    IOPAD_TRI \Q1Q8_pad/U0/U0  (.D(\Q1Q8_pad/U0/NET1 ), .E(
        \Q1Q8_pad/U0/NET2 ), .PAD(Q1Q8));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_17  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m38 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[0] )
        );
    NOR2 
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa_0_a2_0_0  
        (.A(\top_code_0_sd_sacq_choice[3] ), .B(
        \top_code_0_sd_sacq_choice[1] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_3_i_a2_1 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[9]_net_1 ));
    MX2 \scalestate_0/strippluse_RNO_0[11]  (.A(
        \scalestate_0/strippluse_6[11] ), .B(
        \scalestate_0_strippluse[11] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_570 ));
    DFN1E1 \plusestate_0/timecount_1[13]  (.D(
        \plusestate_0/timecount_5[13] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[13] ));
    DFN1 \top_code_0/relay_on[0]  (.D(
        \top_code_0/relay_on_RNO[0]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[0] ));
    AO1 \scalestate_0/timecount_ret_84_RNO  (.A(
        \scalestate_0/OPENTIME[11]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[11] ), .Y(
        \scalestate_0/timecount_20_iv_2[11] ));
    XO1 \bridge_div_0/dataall_RNIEUFH1[2]  (.A(
        \bridge_div_0/count[2]_net_1 ), .B(
        \bridge_div_0/dataall[2]_net_1 ), .C(
        \bridge_div_0/un1_count_1_0[0] ), .Y(
        \bridge_div_0/un1_count_NE_1[0] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n10 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        );
    DFN1E1 \scalestate_0/S_DUMPTIME[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[11]_net_1 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m144  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_145 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_29_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_134_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_2_Y ));
    OR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I0_un1_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[0]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I0_un1_CO1 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[1]  (.A(
        \s_acq_change_0/s_acqnum_5[1] ), .B(
        \s_acq_change_0_s_acqnum[1] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_71 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m208  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[9] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_209 ));
    XO1 \DUMP_0/dump_coder_0/para5_RNIATB71[6]  (.A(
        \DUMP_0/count_0[6] ), .B(\DUMP_0/dump_coder_0/para5[6]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_1[0] ));
    MX2 \state_1ms_0/timecount_RNO_0[11]  (.A(
        \state_1ms_0/timecount_8[11] ), .B(\state_1ms_0_timecount[11] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_78 ));
    NOR3B \DDS_0/dds_coder_0/i_RNO[1]  (.A(
        \DDS_0/dds_coder_0/N_18_mux ), .B(
        \DDS_0/dds_coder_0/m12_2_net_1 ), .C(\DDS_0/count[2] ), .Y(
        \DDS_0/dds_coder_0/i_RNO[1]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m15  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[17] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_16_0 ));
    DFN1E1 \scalestate_0/CUTTIME90[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[2]_net_1 ));
    NOR2A \syn_md_module_1/syn_md_0/count_RNO_0[2]  (.A(
        \syn_md_module_1/syn_md_0/N_52 ), .B(
        \syn_md_module_1/syn_md_0/N_18 ), .Y(
        \syn_md_module_1/syn_md_0/N_25 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[4]  (.D(\top_code_0_scaledatain[4] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[4]_net_1 ));
    DFN1 \DUMP_0/dump_state_0/cs[5]  (.D(
        \DUMP_0/dump_state_0/cs_RNO_0[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0_on_start ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_20  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_20_Y ));
    DFN1 \timer_top_0/state_switch_0/clk_en_scale  (.D(
        \timer_top_0/state_switch_0/clk_en_scale_0_0_a6_0_a5_net_1 ), 
        .CLK(GLA_net_1), .Q(timer_top_0_clk_en_scale));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIC63I1[20]  (.A(
        \sd_acq_top_0/count[20] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[20]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_19[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_1[0] ));
    IOTRI_OB_EB \relay_on_pad[2]/U0/U1  (.D(\relay_on_c[2] ), .E(VCC), 
        .DOUT(\relay_on_pad[2]/U0/NET1 ), .EOUT(
        \relay_on_pad[2]/U0/NET2 ));
    XA1 \PLUSE_0/qq_timer_1/count_RNO[2]  (.A(
        \PLUSE_0/qq_timer_1/count_c1 ), .B(\PLUSE_0/count_7[2] ), .C(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_1/count_n2 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[7]  (.D(
        \top_code_0_halfdata_0[7] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[7] ));
    NOR2A \scalestate_0/strippluse_RNO_1[5]  (.A(\scalestate_0/N_425 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[5] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[25]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[26]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_310 ));
    DFN1E1 \noisestate_0/acqtime[10]  (.D(\top_code_0_noisedata[10] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[10]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_16  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_3_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_167_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_16_Y ));
    DFN1E1 \scalestate_0/CUTTIME180[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[3]_net_1 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_37_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI03Q6[4]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_4[0] ));
    MX2 \scalestate_0/CS_RNIT5AK[10]  (.A(\scalestate_0/CS[11]_net_1 ), 
        .B(\scalestate_0/CS[10]_net_1 ), .S(timer_top_0_clk_en_scale), 
        .Y(\scalestate_0/N_1225 ));
    AX1C \PLUSE_0/bri_timer_0/count_RNO[2]  (.A(\PLUSE_0/count_8[1] ), 
        .B(\PLUSE_0/count_8[0] ), .C(\PLUSE_0/count_8[2] ), .Y(
        \PLUSE_0/bri_timer_0/count_n2 ));
    OA1C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[2]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[1]_net_1 ), .B(\i_6[1] ), 
        .C(\pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_173 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m155  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_156 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[29]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[30]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_484 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[6]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[6] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[6] ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_40  (.A(
        \timer_top_0/timer_0/N_9 ), .B(
        \timer_top_0/timer_0/timedata[14]_net_1 ), .Y(
        \timer_top_0/timer_0/I_40 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m34  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_27 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_34 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_35 ));
    DFN1E1 \top_code_0/cal_data[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[5] ));
    AND2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_22  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT3_E[5] )
        );
    DFN1E0 \DUMP_0/dump_coder_0/para5[2]  (.D(
        \DUMP_0/dump_coder_0/para5_4[2] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[2]_net_1 ));
    NOR3C \ClockManagement_0/clk_div500_0/un1_count_1_I_51  (.A(
        \ClockManagement_0/clk_div500_0/count[6]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/count[7]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_1_1[0] )
        , .Y(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_pog_array_2[0] )
        );
    DFN1E1 \state_1ms_0/M_DUMPTIME[5]  (.D(
        \top_code_0_state_1ms_data[5] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[5]_net_1 ));
    DFN1 \ClockManagement_0/clk_10k_0/count[5]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[5] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[5]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_111  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_111_Y ));
    NOR2B \scalestate_0/timecount_ret_45_RNO_0  (.A(
        \scalestate_0/CUTTIME180[16]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[16] ));
    IOTRI_OB_EB \interupt_pad/U0/U1  (.D(interupt_c), .E(VCC), .DOUT(
        \interupt_pad/U0/NET1 ), .EOUT(\interupt_pad/U0/NET2 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[6]  (.D(
        \top_code_0_sd_sacq_data[6] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[6]_net_1 ));
    NOR3C \scalestate_0/timecount_RNO_3[20]  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[20]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[20] ));
    RAM512X18 #( .MEMORYFILE("RAM_R2C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R2C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_2_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_2_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_0_net ));
    DFN1E1 \scalestate_0/CUTTIME180[18]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1661 ), .Q(\scalestate_0/CUTTIME180[18]_net_1 )
        );
    NOR2A \DDS_0/dds_state_0/para_RNO_3[31]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[32]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_520 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_5  (.A(
        \timer_top_0/dataout[20] ), .B(
        \timer_top_0/timer_0/timedata[20]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_5_Y ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m201  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_202 ));
    DFN1E1 \scalestate_0/PLUSETIME90[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[7]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m70 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[0] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[0]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[13]  (.D(
        \top_code_0_pd_pluse_data[13] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[13]_net_1 ));
    MX2B \state_1ms_0/reset_out_RNO_0  (.A(state_1ms_0_reset_out), .B(
        \state_1ms_0/CS[1]_net_1 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_154 ));
    DFN1E1 \scalestate_0/PLUSETIME180[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[5]_net_1 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[8]_net_1 ));
    DFN1 \DUMP_0/off_on_timer_0/count[3]  (.D(
        \DUMP_0/off_on_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_2[3] ));
    NOR3C \ClockManagement_0/long_timer_0/count_RNIM49U[11]  (.A(
        \ClockManagement_0/long_timer_0/count[7]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[11]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/count[10]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_4 ));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_33  (.A(
        \ClockManagement_0/clk_10k_0/count[1]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_TMP[0] ), .Y(
        \ClockManagement_0/clk_10k_0/I_33_0 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[9]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[10]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_289 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[6] ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[3] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[3]  (.D(
        \top_code_0_bri_datain[7] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[3] ));
    AO1C \timer_top_0/timer_0/Timer_Cmp_0/AO1C_8  (.A(
        \timer_top_0/dataout[21] ), .B(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_0_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_8_Y ));
    NOR2A \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un1_count_0_I_3  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[0]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_4_0 ));
    OA1B \syn_md_module_1/syn_md_0/count_RNO[0]  (.A(
        \syn_md_module_1/syn_md_0/N_23_1 ), .B(
        \syn_md_module_1/syn_md_0/N_28 ), .C(
        \syn_md_module_1/syn_md_0/N_50 ), .Y(
        \syn_md_module_1/syn_md_0/count_RNO_0[0]_net_1 ));
    NOR2 \PLUSE_0/qq_state_0/cs_RNO_1[2]  (.A(\PLUSE_0/i_9[1] ), .B(
        Q3Q6_c), .Y(\PLUSE_0/qq_state_0/N_88 ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_1  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_5_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_3_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_7_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_1_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[8]  (.D(
        \top_code_0_sd_sacq_data[8] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[8]_net_1 ));
    OR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIK5557[2]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_13[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_12[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE[0] ));
    MX2B \top_code_0/k2_RNO_0  (.A(k2_c), .B(\xa_c[0] ), .S(
        \top_code_0/N_12 ), .Y(\top_code_0/N_806 ));
    NOR2A \scalestate_0/strippluse_RNO_1[10]  (.A(\scalestate_0/N_430 )
        , .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[10] ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[6]  (.D(
        \DUMP_0/dump_coder_0/para2_4[6]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[6]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[1] ));
    DFN1E1 \state_1ms_0/CUTTIME[10]  (.D(
        \top_code_0_state_1ms_data[10] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[10]_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[4]  (
        .D(\s_acq_change_0_s_acqnum[4] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[4]_net_1 )
        );
    NOR2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_1_Y ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI4G8R[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_2[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_3[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_9[0] ));
    NOR3B \scalestate_0/STRIPNUM180_NUM_1_sqmuxa_0_a2  (.A(
        \scalestate_0/N_61 ), .B(\scalestate_0/N_64 ), .C(
        \top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ));
    DFN1 \DDS_0/dds_timer_0/count[3]  (.D(\DDS_0/dds_timer_0/count_n3 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[3] ));
    MX2 \state_1ms_0/timecount_RNO_0[17]  (.A(
        \state_1ms_0/timecount_8[17] ), .B(\state_1ms_0_timecount[17] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_84 ));
    AOI1 \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[5]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[1]_net_1 ), .B(\i_6[1] ), 
        .C(\pd_pluse_top_0/pd_pluse_state_0/cs[5]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_176 ));
    INV \bridge_div_0/clk_4f_reg2_RNO  (.A(
        \bridge_div_0/clk_4f_reg1_net_1 ), .Y(
        \bridge_div_0/clk_4f_reg1_i ));
    OA1C \PLUSE_0/qq_state_1/cs_RNO_0[3]  (.A(
        \PLUSE_0/qq_state_1/cs[3]_net_1 ), .B(\PLUSE_0/i_2[3] ), .C(
        Q4Q5_c), .Y(\PLUSE_0/qq_state_1/N_86 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[8]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c6 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n8 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[6]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_60_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[6] ));
    OR3 \scalestate_0/timecount_ret_69_RNO  (.A(
        \scalestate_0/CUTTIME180_m[15] ), .B(
        \scalestate_0/OPENTIME_m[15] ), .C(
        \scalestate_0/timecount_20_iv_3[15] ), .Y(
        \scalestate_0/timecount_20_iv_7[15] ));
    NOR3B \bridge_div_0/count_RNIEMOM7[0]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[0]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIEMOM7[0]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_5  (.A(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .Y(
        \timer_top_0/timer_0/I_5_2 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m5  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[17] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_6_0 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[13]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[13] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_0[13] ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[2]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m288  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_289 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[3]  (.A(\DDS_0/dds_state_0/N_492 )
        , .B(\DDS_0/dds_state_0/N_491 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[3] ), .Y(
        \DDS_0/dds_state_0/N_157 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[13]  (.A(
        \scalestate_0_timecount[13] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_193 ));
    DFN1E1 \top_code_0/pd_pluse_choice[1]  (.D(\GPMI_0_dataout[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_choice_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_choice[1] ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_7_inst  (.A(
        \scalestate_0/necount_inc_0/Rcout_9_net ), .B(
        \scalestate_0/necount[9]_net_1 ), .Y(
        \scalestate_0/necount1[9] ));
    DFN1E1 \top_code_0/sd_sacq_data[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[7] ));
    DFN1P0 \bridge_div_0/clk_4f_reg2  (.D(\bridge_div_0/clk_4f_reg1_i )
        , .CLK(ddsclkout_c), .PRE(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/clk_4f_reg2_i_0 ));
    DFN1C0 \bridge_div_0/clk_4f/U1  (.D(\bridge_div_0/clk_4f/Y ), .CLK(
        ddsclkout_c), .CLR(bri_dump_sw_0_reset_out_0), .Q(
        \bridge_div_0/clk_4f ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[10]_net_1 ));
    INV \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBUBBLEB  (.A(
        top_code_0_n_rd_en), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_119  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_119_Y ));
    NOR2B \scalestate_0/CS_RNO[7]  (.A(\scalestate_0/N_1222 ), .B(
        top_code_0_scale_rst_4), .Y(\scalestate_0/CS_RNO_1[7] ));
    OR3 \DUMP_0/dump_coder_0/para2_RNIK1AT6[0]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_NE_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_3_NE_6[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_3_NE_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_i[0] ));
    MX2 \s_acq_change_0/s_load_0_0_RNIIKH91  (.A(
        \s_acq_change_0/s_load_5_net_1 ), .B(s_acq_change_0_s_load_0), 
        .S(\top_code_0_change[1] ), .Y(\s_acq_change_0/N_69 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[15]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m44_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[15] ));
    AO1 \scalestate_0/timecount_ret_57_RNO_2  (.A(
        \scalestate_0/CUTTIME180_TEL[0]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[0] ), 
        .Y(\scalestate_0/timecount_20_iv_3[0] ));
    DFN1E1 \scalestate_0/ACQTIME[1]  (.D(\top_code_0_scaledatain_0[1] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[1]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_12_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_12_net ));
    DFN1 \top_code_0/relay_close[2]  (.D(
        \top_code_0/relay_close_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[2] ));
    DFN1E1 \top_code_0/dump_sustain_data[2]  (.D(\GPMI_0_dataout[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dump_sustain_data_1_sqmuxa ), 
        .Q(\top_code_0_dump_sustain_data[2] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIU90P[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_11[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_18  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_18_Y ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[2]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_35_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[2] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI5AT7[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_6[0] ));
    DFN1 \top_code_0/relay_on[3]  (.D(
        \top_code_0/relay_on_RNO[3]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[3] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[9]  (.D(
        \top_code_0_state_1ms_data[9] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[9]_net_1 ));
    AO1A \scalestate_0/timecount_ret_65_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[13]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[13] ), .Y(
        \scalestate_0/timecount_20_iv_0[13] ));
    DFN1E1 \scalestate_0/CUTTIME90[20]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[20]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i18_mux ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[10]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_52_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[10] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_7  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[6] )
        );
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[15]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c14 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n15 ));
    DFN1 \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2  (.D(
        \GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_RNO_net_1 ), .CLK(GLA_net_1), 
        .Q(\GPMI_0/xwe_xzcs2_syn_0/xwe_reg2_net_1 ));
    IOPAD_TRI \relay_on_pad[7]/U0/U0  (.D(\relay_on_pad[7]/U0/NET1 ), 
        .E(\relay_on_pad[7]/U0/NET2 ), .PAD(relay_on[7]));
    IOPAD_BI \xd_pad[6]/U0/U0  (.D(\xd_pad[6]/U0/NET1 ), .E(
        \xd_pad[6]/U0/NET2 ), .Y(\xd_pad[6]/U0/NET3 ), .PAD(xd[6]));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[7]  (.A(
        \plusestate_0_timecount[7] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_209 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[12]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[12] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[12] ));
    AO1A \scalestate_0/timecount_ret_23_RNO_0  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[10]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[10] ), .Y(
        \scalestate_0/timecount_20_iv_0[10] ));
    DFN1E1 \scanstate_0/timecount_1[8]  (.D(
        \scanstate_0/timecount_5[8] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[8] ));
    NOR2B \DDS_0/dds_state_0/fq_ud_RNO  (.A(
        \DDS_0/dds_state_0/fq_ud_reg_net_1 ), .B(
        \DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/fq_ud_RNO_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_140  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_14_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_147_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_140_Y ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/FOR2_8_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_10_net ), 
        .B(\pd_pluse_top_0/count_0[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[10] ));
    AO1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO_1[9]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .B(
        \sd_acq_top_0/i_0[7] ), .C(\sd_acq_top_0/sd_sacq_state_0/cs4 ), 
        .Y(\sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[9] ));
    NOR2A \PLUSE_0/bri_state_0/cs_RNO[0]  (.A(
        \PLUSE_0/bri_state_0/cs[0]_net_1 ), .B(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_9[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[12]_net_1 ), 
        .B(\pd_pluse_top_0/count[12] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_12[0] ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[9]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n9 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ));
    DFN1 \sd_acq_top_0/sd_sacq_coder_0/i[3]  (.D(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[3] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/i_5[3] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para1[3]  (.D(
        \top_code_0_bri_datain[3] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para1[3] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[4]  (.D(
        \DUMP_0/dump_coder_0/para5_4[4] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[4]_net_1 ));
    DFN1E1 \top_code_0/dumpdata[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[11] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[4]_net_1 ));
    NOR2A \bridge_div_0/clk_4f_RNO  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/clk_4f ), .Y(\bridge_div_0/clk_4f_5 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[4]  (.A(\s_acq_change_0/N_74 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[4]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[9]_net_1 ));
    NOR3C \DDS_0/dds_coder_0/i_RNO[3]  (.A(\DDS_0/dds_coder_0/m8_2 ), 
        .B(\DDS_0/dds_coder_0/m8_1 ), .C(\DDS_0/dds_coder_0/N_18_mux ), 
        .Y(\DDS_0/dds_coder_0/i_RNO[3]_net_1 ));
    DFN1 \top_code_0/noise_rst_0_0  (.D(
        \top_code_0/noise_rst_0_0_RNIDOO43_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_noise_rst_0));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m281  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[13] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_282 ));
    DFN1E1 \scalestate_0/NE_NUM[2]  (.D(\top_code_0_scaledatain[2] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[2]_net_1 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_42  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[7] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[9] ), .Y(
        \timer_top_0/timer_0/N_8 ));
    IOPAD_TRI \Q4Q5_pad/U0/U0  (.D(\Q4Q5_pad/U0/NET1 ), .E(
        \Q4Q5_pad/U0/NET2 ), .PAD(Q4Q5));
    XO1 \CAL_0/cal_div_0/count_RNII3U71[1]  (.A(
        \CAL_0/cal_para_out[1] ), .B(\CAL_0/cal_div_0/count[1]_net_1 ), 
        .C(\CAL_0/cal_div_0/clear_n4_0 ), .Y(
        \CAL_0/cal_div_0/clear_n4_NE_2 ));
    OR2A \scalestate_0/CS_RNI25262[18]  (.A(\scalestate_0/N_1196 ), .B(
        \scalestate_0/N_1310 ), .Y(\scalestate_0/N_1187 ));
    NOR2B \scalestate_0/CS_RNO[3]  (.A(\scalestate_0/N_1218 ), .B(
        top_code_0_scale_rst_3), .Y(\scalestate_0/CS_RNO_1[3] ));
    DFN1 \timer_top_0/state_switch_0/dataout[18]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[18]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[18] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_54_i ));
    DFN1 \scalestate_0/dumpoff_ctr  (.D(
        \scalestate_0/dumpoff_ctr_RNO_2 ), .CLK(GLA_net_1), .Q(
        scalestate_0_dumpoff_ctr));
    MX2A \scalestate_0/intertodsp_RNO_0  (.A(\scalestate_0/N_1269 ), 
        .B(calcuinter_c), .S(\scalestate_0/un1_CS6_14 ), .Y(
        \scalestate_0/N_727 ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_2  (.A(\ADC_c[8] ), 
        .B(top_code_0_n_s_ctrl_1), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[9]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[9] ));
    OR2A \bri_dump_sw_0/turn_delay_RNO  (.A(top_code_0_pluse_scale), 
        .B(scalestate_0_ne_le), .Y(\bri_dump_sw_0/turn_delay_4 ));
    IOIN_IB \xa_pad[14]/U0/U1  (.YIN(\xa_pad[14]/U0/NET1 ), .Y(
        \xa_c[14] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[7]  (.A(
        \top_code_0_s_acqnum_2[7] ), .B(\scalestate_0_s_acqnum[7] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[7] ));
    IOPAD_IN \XRD_pad/U0/U0  (.PAD(XRD), .Y(\XRD_pad/U0/NET1 ));
    MX2 \state_1ms_0/timecount_RNO_0[15]  (.A(
        \state_1ms_0/timecount_8[15] ), .B(\state_1ms_0_timecount[15] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_82 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/FND2_9_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_12_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_10_net ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_10_net ));
    AO1 \scalestate_0/timecount_ret_14_RNO_2  (.A(
        \scalestate_0/CUTTIME180[9]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[9] ), .Y(
        \scalestate_0/timecount_20_iv_2[9] ));
    XOR2 \PLUSE_0/qq_coder_0/i_reg10_2[0]  (.A(\PLUSE_0/qq_para3[2] ), 
        .B(\PLUSE_0/count_9[2] ), .Y(
        \PLUSE_0/qq_coder_0/i_reg10_2[0]_net_1 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m43  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_38_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m43_5 ));
    DFN1E1 \top_code_0/dump_sustain_data[1]  (.D(\GPMI_0_dataout[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dump_sustain_data_1_sqmuxa ), 
        .Q(\top_code_0_dump_sustain_data[1] ));
    DFN1E1 \scalestate_0/timecount_ret_91  (.D(
        \scalestate_0/timecount_20_iv_6[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[8] ));
    OR3 \scalestate_0/timecount_ret_60_RNIA7I  (.A(
        \scalestate_0/timecount_20_iv_7_reto[12] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[12] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[12] ), .Y(
        \scalestate_0_timecount[12] ));
    NOR2B \state_1ms_0/timecount_RNO_1[19]  (.A(
        \state_1ms_0/CUTTIME[19]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/timecount_8[19] ));
    NOR2 \noisestate_0/CS_RNI1LV7[6]  (.A(\noisestate_0/CS[6]_net_1 ), 
        .B(\noisestate_0/CS[7]_net_1 ), .Y(\noisestate_0/N_250 ));
    MIN3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m4  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[1] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_2_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i2_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[7]_net_1 ));
    DFN1E1 \top_code_0/n_divnum[3]  (.D(\GPMI_0_dataout[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[3] ));
    NOR2B \scalestate_0/timecount_ret_23_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[10]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[10] ));
    NOR2B \dds_change_0/dds_conf_RNO_3  (.A(plusestate_0_dds_config), 
        .B(\top_code_0_change[1] ), .Y(\dds_change_0/dds_confin3_m ));
    OA1A \DDS_0/dds_state_0/w_clk_reg_RNO  (.A(
        \DDS_0/dds_state_0/N_227 ), .B(\DDS_0/dds_state_0/cs[5]_net_1 )
        , .C(\DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/w_clk_reg_RNO_net_1 ));
    OR2B \scalestate_0/pn_out_RNO_2  (.A(\scalestate_0/N_1153_1 ), .B(
        timer_top_0_clk_en_scale), .Y(\scalestate_0/N_1191 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m236  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_237 ));
    OA1C \sd_acq_top_0/sd_sacq_state_0/cs_RNO[9]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/N_207 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[9]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs_srsts_0_i_0[9] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[9]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_124  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_137_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_7_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_124_Y ));
    DFN1E1 \plusestate_0/timecount_1[12]  (.D(
        \plusestate_0/timecount_5[12] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[12] ));
    OR2 \top_code_0/un1_state_1ms_rst_n117_45_i_o2  (.A(
        \top_code_0/N_152 ), .B(\top_code_0/N_157 ), .Y(
        \top_code_0/N_192 ));
    OR3 \scalestate_0/timecount_ret_62_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[12] ), .B(
        \scalestate_0/OPENTIME_TEL_m[12] ), .C(
        \scalestate_0/timecount_20_iv_4[12] ), .Y(
        \scalestate_0/timecount_20_iv_8[12] ));
    DFN1E1 \scalestate_0/PLUSETIME90[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[4]_net_1 ));
    XOR2 \scalestate_0/M_pulse_RNO_6  (.A(
        \scalestate_0/M_NUM[7]_net_1 ), .B(
        \scalestate_0/necount[7]_net_1 ), .Y(\scalestate_0/M_pulse8_7 )
        );
    DFN1E1 \scanstate_0/dectime[4]  (.D(\top_code_0_scandata[4] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[4]_net_1 ));
    NOR2 \noisestate_0/n_acq_RNO_1  (.A(\noisestate_0/CS[4]_net_1 ), 
        .B(\noisestate_0/CS[5]_net_1 ), .Y(\noisestate_0/N_229 ));
    AND3B \DDS_0/dds_coder_0/m3_e  (.A(\DDS_0/count[7] ), .B(
        \DDS_0/count[4] ), .C(\DDS_0/dds_coder_0/m3_e_1_net_1 ), .Y(
        \DDS_0/dds_coder_0/N_18_mux ));
    AO1A \top_code_0/scan_start_ret_3_RNO  (.A(\top_code_0/N_171 ), .B(
        \top_code_0/un1_state_1ms_rst_n117_47_i_a2_0 ), .C(
        \top_code_0/N_162 ), .Y(\top_code_0/N_108 ));
    NOR3B \ClockManagement_0/long_timer_0/timeup_RNO_1  (.A(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_0 ), .B(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_7 ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_7 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_12 ));
    AX1C \PLUSE_0/bri_timer_0/count_RNO[4]  (.A(\PLUSE_0/count_8[3] ), 
        .B(\PLUSE_0/bri_timer_0/count_c2 ), .C(\PLUSE_0/count_8[4] ), 
        .Y(\PLUSE_0/bri_timer_0/count_n4 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[7]  (.A(\scalestate_0/N_455 ), 
        .B(\scalestate_0/ACQECHO_NUM[7]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[7] ));
    DFN1 \DDS_0/dds_timer_0/count[0]  (.D(\DDS_0/dds_timer_0/count_n0 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[0] ));
    AO1 \DDS_0/dds_state_0/para_RNO[0]  (.A(
        \DDS_0/dds_state_0/para[0]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569_0 ), .C(\DDS_0/dds_state_0/N_528 ), 
        .Y(\DDS_0/dds_state_0/N_203 ));
    MX2 \noisestate_0/timecount_1_RNO_0[8]  (.A(
        \noisestate_0/acqtime[8]_net_1 ), .B(
        \noisestate_0/dectime[8]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_65 ));
    DFN1E1 \bridge_div_0/datahalf[1]  (.D(\top_code_0_scaleddsdiv[1] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/datahalf[1]_net_1 ));
    AO1A \state_1ms_0/timecount_RNO_4[2]  (.A(
        \state_1ms_0/S_DUMPTIME[2]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CUTTIME_i_m[2] ), 
        .Y(\state_1ms_0/timecount_8_iv_2[2] ));
    DFN1E1 \state_1ms_0/CUTTIME[13]  (.D(
        \top_code_0_state_1ms_data[13] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[13]_net_1 ));
    DFN1 \plusestate_0/state_over_n  (.D(
        \plusestate_0/state_over_n_RNO_0 ), .CLK(GLA_net_1), .Q(
        plusestate_0_state_over_n));
    NOR2B \scalestate_0/timecount_ret_77_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[6]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[6] ));
    NOR2 \PLUSE_0/qq_state_0/cs_RNO_1[3]  (.A(\PLUSE_0/i_4[2] ), .B(
        \PLUSE_0/qq_state_0/cs[3]_net_1 ), .Y(
        \PLUSE_0/qq_state_0/N_87 ));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_35  (.A(
        \ClockManagement_0/clk_10k_0/count[2]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_1[0] ), .Y(
        \ClockManagement_0/clk_10k_0/I_35_0 ));
    DFN1E1 \noisestate_0/timecount_1[3]  (.D(
        \noisestate_0/timecount_5[3] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[3] ));
    DFN1 \s_acq_change_0/s_stripnum[10]  (.D(
        \s_acq_change_0/s_stripnum_RNO[10]_net_1 ), .CLK(GLA_net_1), 
        .Q(\s_acq_change_0_s_stripnum[10] ));
    NOR3B \timer_top_0/state_switch_0/state_start5_0_0_a2_3  (.A(
        \timer_top_0/state_switch_0/N_285 ), .B(
        \timer_top_0/state_switch_0/N_293 ), .C(
        top_code_0_state_1ms_start), .Y(
        \timer_top_0/state_switch_0/N_297 ));
    NOR2A \scalestate_0/strippluse_RNO_1[1]  (.A(\scalestate_0/N_421 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[1] ));
    NOR2B \DUMP_0/dump_coder_0/para5_RNO[8]  (.A(
        \top_code_0_dumpdata_0[8] ), .B(
        \DUMP_0/dump_coder_0/para19_net_1 ), .Y(
        \DUMP_0/dump_coder_0/para5_4[8] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_62_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIAM0P[17]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[17]_net_1 ), .B(
        \sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_17[0] ));
    AND3 \bridge_div_0/count_5_I_13  (.A(
        \bridge_div_0/DWACT_FINC_E[0] ), .B(
        \bridge_div_0/count_RNIHPOM7[3]_net_1 ), .C(
        \bridge_div_0/count_RNIIQOM7[4]_net_1 ), .Y(\bridge_div_0/N_2 )
        );
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m167  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_168 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m299  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[12] ), .C(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_300 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[8] ));
    DFN1E0 \DDS_0/dds_state_0/para[2]  (.D(\DDS_0/dds_state_0/N_155 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[2]_net_1 ));
    NOR3B \top_code_0/un1_state_1ms_rst_n117_28_i_a2  (.A(
        \top_code_0/N_169 ), .B(\top_code_0/N_334 ), .C(
        \top_code_0/N_152 ), .Y(\top_code_0/N_320 ));
    MX2 \scalestate_0/CS_RNO_0[6]  (.A(\scalestate_0/CS[6]_net_1 ), .B(
        \scalestate_0/CS[5]_net_1 ), .S(timer_top_0_clk_en_scale_0), 
        .Y(\scalestate_0/N_1221 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[3]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[3] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[7]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[7] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_1[7] ));
    NOR2 \top_code_0/relay_close_1_sqmuxa_0_a2_0  (.A(\xa_c[5] ), .B(
        \xa_c[7] ), .Y(\top_code_0/N_337 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[8]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[7] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c6 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n8 ));
    NOR2B \plusestate_0/soft_d_RNO  (.A(\plusestate_0/N_121 ), .B(
        top_code_0_pluse_rst), .Y(\plusestate_0/soft_d_RNO_1_net_1 ));
    IOBI_IB_OB_EB \xd_pad[1]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[1] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[1]/U0/NET3 ), .DOUT(\xd_pad[1]/U0/NET1 ), .EOUT(
        \xd_pad[1]/U0/NET2 ), .Y(\xd_in[1] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIO4QC1[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_4[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_15[0] ));
    AO1A \scalestate_0/timecount_20_iv_4[5]  (.A(\scalestate_0/N_1069 )
        , .B(\scalestate_0/CUTTIME90[5]_net_1 ), .C(
        \scalestate_0/CUTTIMEI90_m[5] ), .Y(
        \scalestate_0/timecount_20_iv_4[5]_net_1 ));
    NOR2A \top_code_0/un1_xa_2_0_a2_0  (.A(\xa_c[4] ), .B(
        \top_code_0/N_158 ), .Y(\top_code_0/N_334 ));
    DFN1E1 \plusestate_0/DUMPTIME[5]  (.D(\top_code_0_plusedata[5] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[5]_net_1 ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[6]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[6]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_2[6] ));
    NOR3B \DUMP_0/off_on_state_0/cs_RNO[1]  (.A(
        state1ms_choice_0_reset_out), .B(\DUMP_0/i_1[0] ), .C(
        \DUMP_0/off_on_state_0/N_10 ), .Y(
        \DUMP_0/off_on_state_0/cs_nsss[1] ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m42_2 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_27[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[3]_net_1 ), .B(
        \sd_acq_top_0/count_10[3] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_3[0] ));
    DFN1 \scalestate_0/strippluse[7]  (.D(
        \scalestate_0/strippluse_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[7] ));
    DFN1E1 \top_code_0/sigtimedata[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[13] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[7]  (.A(
        \scanstate_0_timecount[7] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_206 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m138  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[19] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_139 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m47 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIB6DO6[2]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_9[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_8[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19[0]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_14[0] ));
    NOR3C \timer_top_0/state_switch_0/state_start5_0_0_a2  (.A(
        \timer_top_0/state_switch_0/N_285 ), .B(
        top_code_0_state_1ms_start), .C(
        \timer_top_0/state_switch_0/N_282 ), .Y(
        \timer_top_0/state_switch_0/N_289 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_156  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_156_Y ));
    NOR3C \CAL_0/cal_div_0/count_RNO[2]  (.A(net_33_0), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(\CAL_0/cal_div_0/I_7 ), 
        .Y(\CAL_0/cal_div_0/count_5[2] ));
    NOR2B \DUMP_ON_0/off_on_timer_0/count_RNI96OD[1]  (.A(
        \DUMP_ON_0/count_5[0] ), .B(\DUMP_ON_0/count_5[1] ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_c1 ));
    DFN1E1 \top_code_0/bridge_load  (.D(\top_code_0/N_62 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_bridge_load));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[1] ));
    XOR2 \scalestate_0/necount_inc_0/XOR2_2_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount[3]_net_1 ), .Y(
        \scalestate_0/necount1[3] ));
    NOR2A \syn_md_module_1/syn_md_0/count_RNO_0[0]  (.A(
        \syn_md_module_1/syn_md_0/N_52 ), .B(
        \syn_md_module_1/syn_md_0/count[0]_net_1 ), .Y(
        \syn_md_module_1/syn_md_0/N_28 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[10]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_14_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_4_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_14_net ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[7]  (.D(
        \top_code_0_state_1ms_data[7] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[7]_net_1 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[2]  (.A(\s_acq_change_0/N_58 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[2]_net_1 ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[10]  (.D(
        \top_code_0_state_1ms_data[10] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[10]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[7] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_1  (.A(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .B(
        \timer_top_0/dataout[8] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_1_Y ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNI9ULS[10]  (.A(
        \DUMP_0/dump_coder_0/para2[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_10[0] ));
    NOR3C \DDS_0/dds_timer_0/count_RNO_0[7]  (.A(\DDS_0/count[5] ), .B(
        \DDS_0/dds_timer_0/count_c4 ), .C(
        \DDS_0/dds_timer_0/count_15_0 ), .Y(\DDS_0/dds_timer_0/N_36 ));
    DFN1E1 \top_code_0/scanchoice  (.D(\top_code_0/N_98 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_scanchoice));
    AND3 \timer_top_0/timer_0/un2_timedata_I_48  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[10] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[11] ), .Y(
        \timer_top_0/timer_0/N_6 ));
    DFN1E1 \scalestate_0/timecount_ret_51  (.D(
        \scalestate_0/timecount_20_0_iv_0[18] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_0_reto[18] ));
    DFN1 \PLUSE_0/qq_coder_1/i[1]  (.D(\PLUSE_0/qq_coder_1/i_RNO_7[1] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_7[1] ));
    DFN1E1 \noisestate_0/timecount_1[15]  (.D(
        \noisestate_0/timecount_5[15] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[15] ));
    AND3C \top_code_0/un1_state_1ms_rst_n117_43_i_a3  (.A(\xa_c[4] ), 
        .B(\top_code_0/N_165 ), .C(\top_code_0/N_171 ), .Y(
        \top_code_0/N_327 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/signal_data_t_0_12  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] ), .Y(
        \Signal_Noise_Acq_0/un1_signal_acq_0[2] ));
    IOIN_IB \ADC_pad[0]/U0/U1  (.YIN(\ADC_pad[0]/U0/NET1 ), .Y(
        \ADC_c[0] ));
    OR2 OR2_1 (.A(nsctrl_choice_0_dumpon_ctr), .B(net_40), .Y(OR2_1_Y));
    DFN1E1 \noisestate_0/dectime[5]  (.D(\top_code_0_noisedata[5] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[5]_net_1 ));
    IOBI_IB_OB_EB \xd_pad[13]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[13] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[13]/U0/NET3 ), .DOUT(
        \xd_pad[13]/U0/NET1 ), .EOUT(\xd_pad[13]/U0/NET2 ), .Y(
        \xd_in[13] ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIFM6B5[13]  (.A(
        \ClockManagement_0/long_timer_0/count_c12 ), .B(
        \ClockManagement_0/long_timer_0/count[13]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c13 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[18]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[18] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[18] ));
    DFN1 \noisestate_0/CS[7]  (.D(\noisestate_0/CS_RNO[7]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[7]_net_1 ));
    DFN1E1 \scanstate_0/acqtime[15]  (.D(\top_code_0_scandata[15] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[15]_net_1 ));
    DFN1E1 \top_code_0/state_1ms_data[6]  (.D(\GPMI_0_dataout[6] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[6] ));
    DFN1 \timer_top_0/timer_0/time_up  (.D(
        \timer_top_0/timer_0/time_up_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0_time_up ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m39  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_38_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[16] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_40_i ));
    AX1C \CAL_0/cal_div_0/un3_count_I_7  (.A(
        \CAL_0/cal_div_0/count[1]_net_1 ), .B(
        \CAL_0/cal_div_0/count[0]_net_1 ), .C(
        \CAL_0/cal_div_0/count[2]_net_1 ), .Y(\CAL_0/cal_div_0/I_7 ));
    DFN1 \timer_top_0/state_switch_0/dataout[13]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[13]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[13] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i20_mux ));
    AOI1 \sd_acq_top_0/sd_sacq_state_0/cs_RNO_0[6]  (.A(
        \sd_acq_top_0/i_5[2] ), .B(
        \sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/cs[6]_net_1 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_218 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIS1KG[11]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[11]_net_1 ), .B(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_11[0] ));
    AO1B \scanstate_0/CS_RNO_0[1]  (.A(\scanstate_0/CS_li[0] ), .B(
        timer_top_0_clk_en_scan), .C(net_33_0), .Y(
        \scanstate_0/CS_srsts_i_0[1] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[3]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[3]_net_1 ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_7  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[1]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[2]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_7_1 ));
    DFN1E1 \noisestate_0/dectime[15]  (.D(\top_code_0_noisedata[15] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[15]_net_1 ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNICRST[3]  (
        .A(\pd_pluse_top_0/count_6[3] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[3]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_0[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_7[0] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[3]  (.A(
        \top_code_0_s_acqnum_2[3] ), .B(\scalestate_0_s_acqnum[3] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[3] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI7CT7[7]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[7]_net_1 ), .B(
        \sd_acq_top_0/count_3[7] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_7[0] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[5]  (.D(
        \DUMP_0/dump_coder_0/para5_4[5] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[5]_net_1 ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[9]  (.A(\s_acq_change_0/N_65 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[9]_net_1 ));
    AO1 \scalestate_0/timecount_ret_45_RNO  (.A(
        \scalestate_0/OPENTIME[16]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[16] ), .Y(
        \scalestate_0/timecount_20_0_iv_0[16] ));
    OR2A \scalestate_0/necount_LE_NE_RNI45HP  (.A(top_code_0_scale_rst)
        , .B(\scalestate_0/N_1267 ), .Y(\scalestate_0/N_1206 ));
    DFN1E1 \plusestate_0/DUMPTIME[14]  (.D(\top_code_0_plusedata[14] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[14]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME90[21]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[21]_net_1 ));
    DFN1 \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg2_net_1 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_1_7_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_2_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_5_net ), .C(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_7_net ));
    DFN1 \state_1ms_0/timecount[2]  (.D(
        \state_1ms_0/timecount_RNO[2]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[2] ));
    DFN1E1 \scalestate_0/OPENTIME[17]  (.D(\top_code_0_scaledatain[1] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1681 ), .Q(
        \scalestate_0/OPENTIME[17]_net_1 ));
    DFN1E1 \top_code_0/scaledatain[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[1] ));
    DFN1E1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[1]  
        (.D(\top_code_0_s_periodnum[1] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[1]_net_1 )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[5] ));
    NOR2B \scalestate_0/strippluse_RNO[4]  (.A(\scalestate_0/N_563 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[4]_net_1 ));
    DFN1E1 \top_code_0/halfdata[0]  (.D(\GPMI_0_dataout_0[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[0] ));
    DFN1 \timer_top_0/timer_0/timedata[4]  (.D(
        \timer_top_0/timer_0/timedata_4[4] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[4]_net_1 ));
    AO1A \scalestate_0/timecount_ret_2_RNO_5  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[6]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[6] ), .Y(
        \scalestate_0/timecount_20_iv_1[6] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIU6EN[10]  (.A(
        \sd_acq_top_0/count_1[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[10]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_6[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_5[0] ));
    DFN1 \scalestate_0/s_acqnum_1[9]  (.D(
        \scalestate_0/s_acqnum_1_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_s_acqnum[9] ));
    XA1C \PLUSE_0/qq_coder_0/i_RNO_4[1]  (.A(\PLUSE_0/count_9[3] ), .B(
        \PLUSE_0/qq_para1[3] ), .C(\PLUSE_0/count_9[4] ), .Y(
        \PLUSE_0/qq_coder_0/i_0_0[1] ));
    AO1C \plusestate_0/timecount_1_RNO_1[2]  (.A(
        \plusestate_0/CS[3]_net_1 ), .B(\plusestate_0/N_303 ), .C(
        top_code_0_pluse_rst_0), .Y(\plusestate_0/N_247 ));
    NOR2A \ClockManagement_0/long_timer_0/clk_5K_reg2_RNILRGJ  (.A(
        \ClockManagement_0/long_timer_0/clk_5K_reg1_net_1 ), .B(
        \ClockManagement_0/long_timer_0/clk_5K_reg2_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/clk_5K_en_1 ));
    OR3 \top_code_0/scanchoice_RNO_0  (.A(\top_code_0/N_151 ), .B(
        \top_code_0/N_158 ), .C(\top_code_0/N_157 ), .Y(
        \top_code_0/N_208 ));
    DFN1E1 \top_code_0/pd_pluse_data[5]  (.D(\GPMI_0_dataout[5] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[5] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n4 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[4]_net_1 )
        );
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m45_6 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[7]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[7] ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I9_CO1  
        (.A(\s_acq_change_0_s_stripnum[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N160 ), .C(
        \s_acq_change_0_s_stripnum[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N168 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m256  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_253 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_256 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_257 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[11]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n11 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[11] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m51  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[10] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i18_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_52_i ));
    OR3 \state_1ms_0/timecount_RNO_1[6]  (.A(
        \state_1ms_0/timecount_8_iv_1[6] ), .B(
        \state_1ms_0/timecount_8_iv_0[6] ), .C(
        \state_1ms_0/timecount_8_iv_2[6] ), .Y(
        \state_1ms_0/timecount_8_iv[6] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I5_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I4_un1_CO1 ), 
        .B(\s_acq_change_0_s_stripnum[5] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N152 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_3  
        (.A(\s_acq_change_0_s_stripnum[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N160 ), .C(
        \s_acq_change_0_s_stripnum[9] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_9_0 )
        );
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/ADD_20x20_slow_I19_Y_4 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[19] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m47_3 ));
    AND2 \scalestate_0/necount_inc_0/FND2_8_inst  (.A(
        \scalestate_0/necount_inc_0/incb_2_net ), .B(
        \scalestate_0/necount[9]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/inc_12_net ));
    DFN1E1 \scalestate_0/CUTTIMEI90[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[6]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m102  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_103 ));
    NOR2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y ));
    NOR2B \scalestate_0/timecount_ret_5_RNO_3  (.A(
        \scalestate_0/OPENTIME[2]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[2] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[5]  (.A(\scalestate_0/N_453 ), 
        .B(\scalestate_0/ACQECHO_NUM[5]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[5] ));
    MX2 \nsctrl_choice_0/soft_d_RNO_0  (.A(scanstate_0_soft_d), .B(
        noisestate_0_soft_d), .S(top_code_0_n_s_ctrl_0), .Y(
        \nsctrl_choice_0/soft_d_5 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_37_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_39_i ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIR33A[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[0]_net_1 ), .B(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_0_0[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m164  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_163 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_164 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_165 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_66_i ));
    IOPAD_TRI \Q2Q7_pad/U0/U0  (.D(\Q2Q7_pad/U0/NET1 ), .E(
        \Q2Q7_pad/U0/NET2 ), .PAD(Q2Q7));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[10]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_179 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_180 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[10]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m65  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_66_i ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_7[10]  (.A(
        \sd_acq_top_0/count[16] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[16]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_19[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_2[10] ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[3]_net_1 ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_7  (.A(\ADC_c[3] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_7 ));
    OR3 \scalestate_0/timecount_ret_20_RNIIGA1  (.A(
        \scalestate_0/timecount_20_iv_9_reto[8] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[8] ), .C(
        \scalestate_0/timecount_11_sqmuxa_m_reto ), .Y(
        \scalestate_0_timecount[8] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n1 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[1]_net_1 )
        );
    DFN1E1 \scalestate_0/OPENTIME_TEL[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[15]_net_1 ));
    DFN1 \s_acq_change_0/s_acqnum[4]  (.D(
        \s_acq_change_0/s_acqnum_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[4] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_18[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[7]_net_1 ), .B(
        \pd_pluse_top_0/count_1[7] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_7[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[22]  (.A(
        \DDS_0/dds_state_0/N_538 ), .B(
        \DDS_0/dds_state_0/para[22]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_459 ));
    NOR2B \state_1ms_0/timecount_RNO_5[0]  (.A(
        \state_1ms_0/PLUSECYCLE[0]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[0] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIOSP21[16]  (.A(
        \sd_acq_top_0/count[16] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[16]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_18[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_2[0] ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[9]  (.A(\scalestate_0/N_556 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[9]_net_1 ));
    NOR3A \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_1  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_5_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1C_7_Y ), .C(
        \timer_top_0/dataout[6] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_1_Y ));
    DFN1E1 \scalestate_0/ACQTIME[11]  (.D(\top_code_0_scaledatain[11] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[11]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_64_i ));
    MX2 \scalestate_0/bb_ch_RNO_0  (.A(\scalestate_0/N_297 ), .B(
        net_51), .S(\scalestate_0/N_1177 ), .Y(\scalestate_0/N_729 ));
    NOR2B \scalestate_0/timecount_ret_87_RNO_0  (.A(
        \scalestate_0/CUTTIME180[10]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[10] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[1]  (.A(
        \scalestate_0_timecount[1] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_238 ));
    NOR3C \DUMP_0/off_on_timer_0/count_0_sqmuxa  (.A(
        \DUMP_0/off_on_state_0_state_over ), .B(
        \DUMP_0/dump_state_0_off_start ), .C(
        state1ms_choice_0_reset_out), .Y(
        \DUMP_0/off_on_timer_0/count_0_sqmuxa_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[6]  (.A(
        \top_code_0_dumpdata_0[6] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[6]_net_1 ));
    DFN1E1 \scanstate_0/timecount_1[3]  (.D(
        \scanstate_0/timecount_5[3] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[3] ));
    DFN1E1 \scalestate_0/ACQ180_NUM[0]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[0]_net_1 ));
    NOR2B \scalestate_0/pluse_start_RNO  (.A(\scalestate_0/N_725 ), .B(
        top_code_0_scale_rst_3), .Y(
        \scalestate_0/pluse_start_RNO_0_net_1 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m36  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[16] ), .B(
        \top_code_0_s_addchoice_4[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_37 ));
    NOR3A \top_code_0/pluse_str_RNO_4  (.A(\xa_c[7] ), .B(
        \top_code_0/N_139 ), .C(\top_code_0/N_190 ), .Y(
        \top_code_0/N_319 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[8]  (
        .D(\s_acq_change_0_s_acqnum[8] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[8]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m158  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_151 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_158 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_159 ));
    AO1 \scalestate_0/timecount_ret_1_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[5]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[5] ), 
        .Y(\scalestate_0/timecount_20_iv_3[5] ));
    NOR3 \top_code_0/sd_sacq_load_RNO_1  (.A(\top_code_0/N_148 ), .B(
        \top_code_0/N_163 ), .C(\top_code_0/N_157 ), .Y(
        \top_code_0/N_310 ));
    NOR2A \plusestate_0/timecount_1_RNO[14]  (.A(\plusestate_0/N_85 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[14] ));
    IOPAD_TRI \relay_on_pad[4]/U0/U0  (.D(\relay_on_pad[4]/U0/NET1 ), 
        .E(\relay_on_pad[4]/U0/NET2 ), .PAD(relay_on[4]));
    XOR2 \CAL_0/cal_div_0/un3_count_I_14  (.A(\CAL_0/cal_div_0/N_2 ), 
        .B(\CAL_0/cal_div_0/count[5]_net_1 ), .Y(
        \CAL_0/cal_div_0/I_14 ));
    DFN1 \dds_change_0/dds_rst  (.D(\dds_change_0/dds_rst_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(dds_change_0_dds_rst));
    MX2 \scanstate_0/timecount_1_RNO_0[1]  (.A(
        \scanstate_0/acqtime[1]_net_1 ), .B(
        \scanstate_0/dectime[1]_net_1 ), .S(\scanstate_0/N_194 ), .Y(
        \scanstate_0/N_59 ));
    OR3 \scalestate_0/timecount_ret_40_RNIJ4EE  (.A(
        \scalestate_0/timecount_20_iv_7_reto[2] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[2] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[2] ), .Y(
        \scalestate_0/timecount_20_iv_10_reto[2] ));
    NOR2B \scalestate_0/CS_RNIRUEO[10]  (.A(\scalestate_0/N_1225 ), .B(
        top_code_0_scale_rst_5), .Y(
        \scalestate_0/CS_RNIRUEO[10]_net_1 ));
    IOPAD_TRI \relay_on_pad[3]/U0/U0  (.D(\relay_on_pad[3]/U0/NET1 ), 
        .E(\relay_on_pad[3]/U0/NET2 ), .PAD(relay_on[3]));
    NOR2 \DDS_0/dds_state_0/cs_RNIB4FB[7]  (.A(
        \DDS_0/dds_state_0/cs[7]_net_1 ), .B(
        \DDS_0/dds_state_0/cs[8]_net_1 ), .Y(\DDS_0/dds_state_0/N_451 )
        );
    DFN1E1 \top_code_0/plusedata[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[1] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m13  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i6_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[4] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i8_mux ));
    NOR2A \ClockManagement_0/clk_10k_0/clk_5M_reg2_RNI337M  (.A(
        \ClockManagement_0/clk_10k_0/clk_5M_reg1_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/clk_5M_reg2_net_1 ), .Y(
        \ClockManagement_0/clk_5M_en ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m43  
        (.A(\s_acq_change_0_s_stripnum[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[10]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i18_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_44_i ));
    DFN1 \ClockManagement_0/clk_10k_0/count[6]  (.D(
        \ClockManagement_0/clk_10k_0/count_5[6] ), .CLK(GLA_net_1), .Q(
        \ClockManagement_0/clk_10k_0/count[6]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[20]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1723 ), .Q(
        \scalestate_0/CUTTIME180_TEL[20]_net_1 ));
    MX2 \PLUSE_0/bri_state_0/down/U0  (.A(\PLUSE_0/down ), .B(
        \PLUSE_0/bri_state_0/down32 ), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_state_0/down/Y ));
    NOR2A \state_1ms_0/CS_i_RNI9BAF[0]  (.A(
        \state_1ms_0/CS_i[0]_net_1 ), .B(\state_1ms_0/CS[9]_net_1 ), 
        .Y(\state_1ms_0/N_257 ));
    XA1 \DUMP_0/off_on_timer_1/count_RNO[3]  (.A(
        \DUMP_0/off_on_timer_1/count_c2 ), .B(\DUMP_0/count_0[3] ), .C(
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_1/count_n3 ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6_RNO_0  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I6_un1_CO1 ), 
        .B(\s_acq_change_0_s_stripnum[7] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_7 ));
    NOR3C \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_2_i ));
    MX2B \topctrlchange_0/interupt_RNO_0  (.A(interupt_c), .B(
        \topctrlchange_0/un1_interin1[0] ), .S(
        \dds_change_0.un1_change_2 ), .Y(\topctrlchange_0/N_8 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m294  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_287 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_294 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[13] ));
    NOR3A \sd_acq_top_0/sd_sacq_state_0/cs_RNO[6]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs4 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/N_218 ), .C(
        \sd_acq_top_0/sd_sacq_state_0/N_219 ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_2[6] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI8M0I[1]  (.A(
        \sd_acq_top_0/count_10[1] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[1]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_9[0] ));
    AO1 \scalestate_0/timecount_ret_68_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[14]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[14] ), .Y(
        \scalestate_0/timecount_20_iv_4[14] ));
    DFN1E1 \scalestate_0/CUTTIME90[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[1]_net_1 ));
    NOR2B \DDS_0/dds_state_0/para_reg_100_e_1  (.A(
        top_code_0_dds_choice), .B(top_code_0_dds_load), .Y(
        \DDS_0/dds_state_0/N_569_1 ));
    DFN1E1 \plusestate_0/DUMPTIME[6]  (.D(\top_code_0_plusedata[6] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[6]_net_1 ));
    NOR3A \sd_acq_top_0/sd_sacq_coder_0/i_RNO_12[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_10[10] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_15[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_1[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_16[10] ));
    AO1B \noisestate_0/state_over_n_RNO  (.A(noisestate_0_state_over_n)
        , .B(\noisestate_0/N_250 ), .C(top_code_0_noise_rst_0), .Y(
        \noisestate_0/state_over_n_RNO_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[13]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_nsss[13] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[13]_net_1 ));
    DFN1 \DUMP_OFF_1/off_on_timer_0/count[4]  (.D(
        \DUMP_OFF_1/off_on_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_1/count_4[4] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_50_i ));
    DFN1E1 \scalestate_0/DUMPTIME[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[15]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[7] ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ));
    DFN1C0 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11]/U1  (
        .D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] ));
    DFN1E0 \DDS_0/dds_state_0/para[14]  (.D(\DDS_0/dds_state_0/N_121 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1_0 ), .Q(
        \DDS_0/dds_state_0/para[14]_net_1 ));
    NOR2B \state_1ms_0/timecount_RNO[1]  (.A(\state_1ms_0/N_68 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/timecount_RNO[1]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[3]_net_1 ));
    DFN1 \DUMP_0/off_on_timer_0/count[0]  (.D(
        \DUMP_0/off_on_timer_0/count_n0 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_2[0] ));
    NAND3A \scalestate_0/necount_cmp_0/NAND3A_2  (.A(
        \scalestate_0/M_NUM[4]_net_1 ), .B(
        \scalestate_0/necount[4]_net_1 ), .C(
        \scalestate_0/necount_cmp_0/OR2A_0_Y ), .Y(
        \scalestate_0/necount_cmp_0/NAND3A_2_Y ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[6]  (.A(
        \timer_top_0/state_switch_0/N_212 ), .B(
        \timer_top_0/state_switch_0/N_214 ), .C(
        \timer_top_0/state_switch_0/N_213 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[6] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_13  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[15]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ADD_16x16_slow_I15_Y )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[2] )
        );
    NOR3C \timer_top_0/timer_0/timedata_RNO[13]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_37_1 ), .Y(
        \timer_top_0/timer_0/timedata_4[13] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNIU3KG[12]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[12]_net_1 ), .B(
        \sd_acq_top_0/count_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_12[0] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m170  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_171 ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_1  (.A(\ADC_c[9] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[10]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[12]  (.D(
        \top_code_0_scaledatain[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[12]_net_1 )
        );
    NOR3 \DDS_0/dds_state_0/para_RNO[14]  (.A(
        \DDS_0/dds_state_0/N_464 ), .B(\DDS_0/dds_state_0/N_463 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[14] ), .Y(
        \DDS_0/dds_state_0/N_121 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[2]  (.D(
        \ClockManagement_0/long_timer_0/count_n2 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[2]_net_1 ));
    DFN1E1 \scalestate_0/NE_NUM[8]  (.D(\top_code_0_scaledatain[8] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[8]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_67  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_67_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[13]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_69_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[15]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[15] ));
    DFN1E1 \scalestate_0/PLUSETIME90[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[6]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[24]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[25]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_305 ));
    DFN1E1 \top_code_0/s_addchoice_2[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_2[0] ));
    NOR2B \top_code_0/k1_RNO  (.A(\top_code_0/N_807 ), .B(net_27), .Y(
        \top_code_0/k1_RNO_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[0]  (.A(
        \top_code_0_dumpdata_0[0] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[0]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[12]_net_1 ));
    DFN1 \state_1ms_0/timecount[7]  (.D(
        \state_1ms_0/timecount_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[7] ));
    NOR3 \timer_top_0/state_switch_0/state_start5_0_0_a2_5  (.A(
        top_code_0_scan_start), .B(top_code_0_noise_start), .C(
        top_code_0_scale_start), .Y(\timer_top_0/state_switch_0/N_285 )
        );
    NOR2 \top_code_0/un1_state_1ms_rst_n117_43_i_a2_0_0  (.A(
        \top_code_0/N_157 ), .B(\top_code_0/N_144 ), .Y(
        \top_code_0/un1_state_1ms_rst_n117_43_i_a2_0_0_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m182  (.A(
        \top_code_0_s_addchoice_2[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[11] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_183 ));
    DFN1E1 \scalestate_0/STRIPNUM180_NUM[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM180_NUM[8]_net_1 ));
    DFN1 \state_1ms_0/CS[9]  (.D(\state_1ms_0/CS_RNO_1[9] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[9]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_23_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[10]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[10] ));
    NOR2B \dds_change_0/dds_conf_RNO  (.A(\dds_change_0/N_6 ), .B(
        net_27), .Y(\dds_change_0/dds_conf_RNO_net_1 ));
    AO1B \state_1ms_0/timecount_RNO_3[1]  (.A(
        \state_1ms_0/M_DUMPTIME[1]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/CS_i[0]_net_1 ), 
        .Y(\state_1ms_0/timecount_8_iv_0[1] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_123  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_123_Y ));
    NOR3 \DDS_0/dds_state_0/para_RNO[16]  (.A(
        \DDS_0/dds_state_0/N_297 ), .B(\DDS_0/dds_state_0/N_296 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[16] ), .Y(
        \DDS_0/dds_state_0/N_18 ));
    DFN1E1 \top_code_0/n_acqnum[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_acqnum_1_sqmuxa ), .Q(
        \top_code_0_n_acqnum_2[11] ));
    DFN1E1 \top_code_0/halfdata[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[2] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[10]  (.A(
        \state_1ms_0_timecount[10] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_252 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_151  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_2_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_2_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_151_Y ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[0]  (.D(
        \top_code_0_state_1ms_data[0] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[0]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME[0]  (.D(\top_code_0_scaledatain[0] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/N_1665 ), .Q(
        \scalestate_0/OPENTIME[0]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_62  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_62_Y ));
    OR3 \scalestate_0/M_pulse_RNO_1  (.A(\scalestate_0/M_pulse8_NE_4 ), 
        .B(\scalestate_0/M_pulse8_NE_3 ), .C(
        \scalestate_0/M_pulse8_NE_8 ), .Y(\scalestate_0/M_pulse8_NE ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[5]  (.A(\scalestate_0/N_552 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[5]_net_1 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para2[1]  (.D(
        \top_code_0_bri_datain[5] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para2[1] ));
    IOPAD_TRI \interupt_pad/U0/U0  (.D(\interupt_pad/U0/NET1 ), .E(
        \interupt_pad/U0/NET2 ), .PAD(interupt));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[14]  (.A(
        \scanstate_0_timecount[14] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_261 ));
    NOR3C \scalestate_0/timecount_ret_2_RNO_6  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[6]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[6] ));
    NOR2A \scalestate_0/strippluse_RNO_1[7]  (.A(\scalestate_0/N_427 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[7] ));
    IOPAD_BI \xd_pad[7]/U0/U0  (.D(\xd_pad[7]/U0/NET1 ), .E(
        \xd_pad[7]/U0/NET2 ), .Y(\xd_pad[7]/U0/NET3 ), .PAD(xd[7]));
    NOR2B \s_acq_change_0/s_acqnum_RNO[13]  (.A(\s_acq_change_0/N_83 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[13]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIS66B[0]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[0]_net_1 ), .B(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_0_0[0] ));
    DFN1E1 \noisestate_0/timecount_1[14]  (.D(
        \noisestate_0/timecount_5[14] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[14] ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[8]  (.D(
        \DUMP_0/dump_coder_0/para2_4[8]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[8]_net_1 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[9]  (.A(
        \s_acq_change_0/s_acqnum_5[9] ), .B(
        \s_acq_change_0_s_acqnum[9] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_79 ));
    XA1 \DUMP_OFF_1/off_on_timer_0/count_RNO[1]  (.A(
        \DUMP_OFF_1/count_4[1] ), .B(\DUMP_OFF_1/count_4[0] ), .C(
        \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_n1 ));
    NOR2B \state_1ms_0/timecount_RNO_6[4]  (.A(
        \state_1ms_0/PLUSETIME[4]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[4] ));
    MX2A \scalestate_0/dump_start_RNO_0  (.A(\scalestate_0/N_1210 ), 
        .B(scalestate_0_dump_start), .S(\scalestate_0/N_1167 ), .Y(
        \scalestate_0/N_723 ));
    OR3 \top_code_0/dumpload_RNO_0  (.A(\top_code_0/N_144 ), .B(
        \top_code_0/N_148 ), .C(\top_code_0/N_164 ), .Y(
        \top_code_0/N_218 ));
    DFN1 \top_code_0/k1  (.D(\top_code_0/k1_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(k1_c));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[7]  (.D(
        \top_code_0_n_acqnum_2[7] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[7]_net_1 ));
    NOR2B \scalestate_0/dds_conf_RNO  (.A(\scalestate_0/N_728 ), .B(
        top_code_0_scale_rst), .Y(\scalestate_0/dds_conf_RNO_0_net_1 ));
    IOBI_IB_OB_EB \xd_pad[6]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[6] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[6]/U0/NET3 ), .DOUT(\xd_pad[6]/U0/NET1 ), .EOUT(
        \xd_pad[6]/U0/NET2 ), .Y(\xd_in[6] ));
    OR3 \DUMP_0/dump_state_0/off_start_RNO_0  (.A(
        \DUMP_0/dump_state_0/N_196 ), .B(\DUMP_0/dump_state_0/N_195 ), 
        .C(\DUMP_0/dump_state_0/N_171 ), .Y(
        \DUMP_0/dump_state_0/N_176 ));
    DFN1E1 \top_code_0/dds_configdata[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[14] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/m45_1 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[14] ));
    XNOR2 \PLUSE_0/bri_coder_0/half_0_I_3  (.A(\PLUSE_0/half_para[5] ), 
        .B(\PLUSE_0/count_2[5] ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_BL_EQUAL_0_E[0] ));
    DFN1 \top_code_0/relay_on[7]  (.D(
        \top_code_0/relay_on_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[7] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIGMR21[20]  (.A(
        \sd_acq_top_0/count[20] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[20]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_19[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_1[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_94  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_129_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_17_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_94_Y ));
    AO1A \state_1ms_0/timecount_RNO_4[6]  (.A(
        \state_1ms_0/S_DUMPTIME[6]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CUTTIME_i_m[6] ), 
        .Y(\state_1ms_0/timecount_8_iv_2[6] ));
    OR3 \scalestate_0/timecount_ret_35_RNO  (.A(
        \scalestate_0/CUTTIMEI90_m[9] ), .B(
        \scalestate_0/CUTTIME90_m[9] ), .C(
        \scalestate_0/timecount_20_iv_5[9] ), .Y(
        \scalestate_0/timecount_20_iv_8[9] ));
    OR2A \PLUSE_0/bri_coder_0/half_0_I_14  (.A(\PLUSE_0/count_8[1] ), 
        .B(\PLUSE_0/half_para[1] ), .Y(\PLUSE_0/bri_coder_0/N_2 ));
    OR3A \top_code_0/RAM_Rd_rst_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_155 ), .C(\top_code_0/N_165 ), .Y(
        \top_code_0/N_206 ));
    NOR2A \sd_acq_top_0/sd_sacq_state_0/cs_RNIIF5E[7]  (.A(
        \sd_acq_top_0/sd_sacq_state_0/cs[7]_net_1 ), .B(
        \sd_acq_top_0/i_0[6] ), .Y(
        \sd_acq_top_0/sd_sacq_state_0/N_235 ));
    NOR2B \top_code_0/relay_close_RNO[0]  (.A(\top_code_0/N_819 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[0]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[22]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[22]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_460 ));
    DFN1E1 \state_1ms_0/CUTTIME[15]  (.D(
        \top_code_0_state_1ms_data[15] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[15]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m137  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_136 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_137 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_138 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_142  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_49_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_10_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_3_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_142_Y ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[0]_net_1 ));
    DFN1E1 \scalestate_0/M_NUM[2]  (.D(\top_code_0_scaledatain_0[2] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[2]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[3]  (.A(
        \noisestate_0/acqtime[3]_net_1 ), .B(
        \noisestate_0/dectime[3]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_60 ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIBMOK[0]  (.A(
        \DUMP_0/dump_coder_0/para6[0]_net_1 ), .B(\DUMP_0/count_1[0] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_0[0] ));
    NOR2A \Signal_Noise_Acq_0/n_s_change_0/s_adc_1_10  (.A(\ADC_c[0] ), 
        .B(top_code_0_n_s_ctrl), .Y(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ));
    NOR3B \DUMP_OFF_1/off_on_coder_0/i_RNO_1[1]  (.A(
        \DUMP_OFF_1/count_4[4] ), .B(\DUMP_OFF_1/count_4[2] ), .C(
        \DUMP_OFF_1/count_4[3] ), .Y(
        \DUMP_OFF_1/off_on_coder_0/i_0_2[1] ));
    DFN1 \syn_md_module_1/syn_md_0/count[2]  (.D(
        \syn_md_module_1/syn_md_0/count_RNO[2]_net_1 ), .CLK(GLA_net_1)
        , .Q(\syn_md_module_1/syn_md_0/count[2]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[8]  (.D(
        \top_code_0_pd_pluse_data[8] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[8]_net_1 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[3]  (.D(
        \top_code_0_halfdata_0[3] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[3] ));
    AO1B \scalestate_0/CS_RNIR1C72[18]  (.A(\scalestate_0/N_1310 ), .B(
        timer_top_0_clk_en_scale_0), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/un1_CS6_33_0 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[5]  (.A(
        \scalestate_0/ACQ180_NUM[5]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[5]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_453 ));
    MX2 \DSTimer_0/dump_sustain_timer_0/data_RNO_0[1]  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[1]_net_1 ), .B(
        \top_code_0_dump_sustain_data[1] ), .S(\DSTimer_0/AND2_0_Y ), 
        .Y(\DSTimer_0/dump_sustain_timer_0/N_25 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[21]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[21] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[21] ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[9]  (.A(
        \PLUSE_0/bri_state_0/cs[9]_net_1 ), .B(
        \PLUSE_0/bri_state_0/N_145 ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[9] ));
    MX2A \scalestate_0/CS_RNO_0[21]  (.A(\scalestate_0/CS[21]_net_1 ), 
        .B(\scalestate_0/N_1208 ), .S(timer_top_0_clk_en_scale_0), .Y(
        \scalestate_0/N_1236 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[1]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n1 ));
    DFN1E1 \noisestate_0/dectime[2]  (.D(\top_code_0_noisedata[2] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[2]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m293  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_290 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_293 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_294 ));
    DFN1E1 \noisestate_0/dectime[8]  (.D(\top_code_0_noisedata[8] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[8]_net_1 ));
    DFN1E1 \scalestate_0/DUMPTIME[6]  (.D(\top_code_0_scaledatain[6] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[6]_net_1 ));
    OA1B \scanstate_0/CS_RNO[4]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[4]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[4] ), 
        .Y(\scanstate_0/CS_RNO_2[4] ));
    MX2C \DUMP_OFF_0/off_on_state_0/cs_RNO_0[1]  (.A(
        \DUMP_OFF_0/off_on_state_0/cs[1]_net_1 ), .B(
        \DUMP_OFF_0/i_3[1] ), .S(DUMP_OFF_0_dump_off), .Y(
        \DUMP_OFF_0/off_on_state_0/N_10 ));
    AX1C \DDS_0/dds_timer_0/count_RNO[7]  (.A(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .B(\DDS_0/count[7] )
        , .C(\DDS_0/dds_timer_0/N_36 ), .Y(
        \DDS_0/dds_timer_0/count_n7 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_159  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_5_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_5_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_159_Y ));
    IOPAD_IN \xa_pad[6]/U0/U0  (.PAD(xa[6]), .Y(\xa_pad[6]/U0/NET1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[3]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[6]  (.D(\GPMI_0_dataout[6] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[6] ));
    NOR2B \scalestate_0/intertodsp_RNO  (.A(\scalestate_0/N_727 ), .B(
        top_code_0_scale_rst_3), .Y(
        \scalestate_0/intertodsp_RNO_0_net_1 ));
    DFN1E1 \state_1ms_0/CUTTIME[7]  (.D(\top_code_0_state_1ms_data[7] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[7]_net_1 ));
    OR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_6 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_7 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_6_net_1 )
        );
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[1] ));
    DFN1E1 \plusestate_0/timecount_1[10]  (.D(
        \plusestate_0/timecount_5[10] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[10] ));
    RAM512X18 #( .MEMORYFILE("RAM_R13C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R13C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_13_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_13_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_0_net )
        );
    XOR2 \bridge_div_0/dataall_1_I_7  (.A(\top_code_0_scaleddsdiv[1] ), 
        .B(\top_code_0_scaleddsdiv[4] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0[0] ));
    AO1A \top_code_0/inv_turn_RNO_1  (.A(\top_code_0/N_167 ), .B(
        \top_code_0/N_340 ), .C(\top_code_0/N_322 ), .Y(
        \top_code_0/N_122 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[8]  (.D(
        \top_code_0_scaledatain[8] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[8]_net_1 ));
    NOR2B \DUMP_OFF_1/off_on_timer_0/count_RNI761C[1]  (.A(
        \DUMP_OFF_1/count_4[0] ), .B(\DUMP_OFF_1/count_4[1] ), .Y(
        \DUMP_OFF_1/off_on_timer_0/count_c1 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[7]  (.A(
        \ClockManagement_0/long_timer_0/count_c6 ), .B(
        \ClockManagement_0/long_timer_0/count[7]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n7 ));
    IOPAD_IN \ADC_pad[3]/U0/U0  (.PAD(ADC[3]), .Y(\ADC_pad[3]/U0/NET1 )
        );
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[15]  (.D(
        \top_code_0_pd_pluse_data[15] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[15]_net_1 ));
    AND2 \DSTimer_0/AND2_0  (.A(\DSTimer_0/net_0 ), .B(
        \DSTimer_0/DFI0_1_QN ), .Y(\DSTimer_0/AND2_0_Y ));
    OR2B \scanstate_0/CS_RNI97DM[1]  (.A(\scanstate_0/CS[1]_net_1 ), 
        .B(net_33), .Y(\scanstate_0/N_196 ));
    DFN1E1 \scalestate_0/PLUSETIME180[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[15]_net_1 ));
    MIN3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m4  (.A(
        \top_code_0_n_divnum_0[1] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_2_i ), .C(
        \top_code_0_n_divnum_0[6] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i2_mux ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[24]  (.D(
        \top_code_0_dds_configdata[7] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[24]_net_1 ));
    DFN1E1 \top_code_0/n_s_ctrl_1  (.D(\top_code_0/N_76 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_n_s_ctrl_1));
    NOR3C \timer_top_0/timer_0/timedata_RNO[11]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_32_2 ), .Y(
        \timer_top_0/timer_0/timedata_4[11] ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_12_RNO_5  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[1]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_1_0 )
        );
    NOR3A \top_code_0/un1_state_1ms_rst_n117_21_i_a2  (.A(
        \top_code_0/N_169 ), .B(\top_code_0/N_154 ), .C(
        \top_code_0/N_148 ), .Y(\top_code_0/N_321 ));
    OR3 \scalestate_0/timecount_ret_23_RNIRFA1  (.A(
        \scalestate_0/timecount_20_iv_9_reto[10] ), .B(
        \scalestate_0/timecount_20_iv_8_reto[10] ), .C(
        \scalestate_0/timecount_11_sqmuxa_m_reto ), .Y(
        \scalestate_0_timecount[10] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[31]  (.A(
        \DDS_0/dds_state_0/N_518 ), .B(\DDS_0/dds_state_0/N_517 ), .C(
        \DDS_0/dds_state_0/para_9_i_0[31] ), .Y(
        \DDS_0/dds_state_0/N_171 ));
    DFN1 \timer_top_0/timer_0/timedata[8]  (.D(
        \timer_top_0/timer_0/timedata_4[8] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[8]_net_1 ));
    MX2C \DUMP_0/off_on_state_1/cs_RNO_0[1]  (.A(
        \DUMP_0/off_on_state_1/cs[1]_net_1 ), .B(\DUMP_0/i_0[1] ), .S(
        DUMP_0_dump_on), .Y(\DUMP_0/off_on_state_1/N_10 ));
    NOR2B \scalestate_0/long_opentime_RNO  (.A(\scalestate_0/N_743 ), 
        .B(top_code_0_scale_rst_3), .Y(
        \scalestate_0/long_opentime_RNO_net_1 ));
    MX2B \plusestate_0/timecount_1_RNO[4]  (.A(\plusestate_0/N_75 ), 
        .B(\plusestate_0/N_249 ), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[4] ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[3]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[3]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_8[3] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[7]  (.D(
        \top_code_0_pd_pluse_data[7] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[7]_net_1 ));
    AO1 \scalestate_0/timecount_ret_19_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL[8]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[8] ), 
        .Y(\scalestate_0/timecount_20_iv_3[8] ));
    XA1 \PLUSE_0/qq_timer_0/count_RNO[4]  (.A(
        \PLUSE_0/qq_timer_0/count_9_0 ), .B(\PLUSE_0/count_9[4] ), .C(
        \PLUSE_0/qq_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_0/count_n4 ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[4]  (.A(\scalestate_0/N_551 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/s_acqnum_1_RNO[4]_net_1 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[8]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_23_0 ), .Y(
        \timer_top_0/timer_0/timedata_4[8] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[5]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c4 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n5 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[1]  (.A(
        \timer_top_0/state_switch_0/N_237 ), .B(
        \timer_top_0/state_switch_0/N_239 ), .C(
        \timer_top_0/state_switch_0/N_238 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[1] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_2[8]  (.A(
        \scalestate_0/ACQ180_NUM[8]_net_1 ), .B(
        \scalestate_0/ACQ90_NUM[8]_net_1 ), .S(\scalestate_0/N_1209 ), 
        .Y(\scalestate_0/N_456 ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa_0_a2  (
        .A(\top_code_0_sd_sacq_choice[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/N_24 ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ));
    NOR2B \state_1ms_0/timecount_RNO_6[0]  (.A(
        \state_1ms_0/PLUSETIME[0]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[0] ));
    DFN1 \scalestate_0/CS[19]  (.D(\scalestate_0/CS_RNO[19]_net_1 ), 
        .CLK(GLA_net_1), .Q(\scalestate_0/CS[19]_net_1 ));
    MX2 \PLUSE_0/bri_timer_0/count[1]/U0  (.A(\PLUSE_0/count_8[1] ), 
        .B(\PLUSE_0/bri_timer_0/count_n1 ), .S(
        \PLUSE_0/bri_timer_0/clken_net_1 ), .Y(
        \PLUSE_0/bri_timer_0/count[1]/Y ));
    XOR2 \ClockManagement_0/clk_div500_0/un1_count_1_I_34  (.A(
        \ClockManagement_0/clk_div500_0/count[6]_net_1 ), .B(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_11[0] ), 
        .Y(\ClockManagement_0/clk_div500_0/I_34 ));
    NOR2B \DUMP_0/off_on_timer_0/count_RNIH8RC[1]  (.A(
        \DUMP_0/count_2[1] ), .B(\DUMP_0/count_2[0] ), .Y(
        \DUMP_0/off_on_timer_0/count_c1 ));
    DFN1 \s_acq_change_0/s_acqnum[5]  (.D(
        \s_acq_change_0/s_acqnum_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[5] ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[15]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[15] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_0[15] ));
    MX2 \dds_change_0/dds_conf_RNO_0  (.A(dds_change_0_dds_conf), .B(
        \dds_change_0/dds_conf_6 ), .S(\dds_change_0.un1_change_2 ), 
        .Y(\dds_change_0/N_6 ));
    DFN1E1 \top_code_0/dumpdata[10]  (.D(\GPMI_0_dataout[10] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[10] ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_5  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[11] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[11]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[4] )
        );
    DFN1E1 \scalestate_0/NE_NUM[9]  (.D(\top_code_0_scaledatain[9] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/NE_NUM_1_sqmuxa ), .Q(
        \scalestate_0/NE_NUM[9]_net_1 ));
    DFN1E1 \scalestate_0/DUMPTIME[0]  (.D(\top_code_0_scaledatain[0] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[0]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[15]  (.D(
        \top_code_0_pd_pluse_data[15] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[15]_net_1 ));
    OA1B \plusestate_0/CS_RNO[7]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[7]_net_1 ), .C(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Y(
        \plusestate_0/CS_RNO_0[7] ));
    MAJ3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I3_CO1  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/perioddata[3]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I2_un1_CO1 ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N146 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[31]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[31]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_518 ));
    DFN1C0 \PLUSE_0/bri_state_0/cs[14]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO[14]_net_1 ), .CLK(ddsclkout_c), 
        .CLR(\PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs[14]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO[8]  (.A(\noisestate_0/N_65 ), .B(
        \noisestate_0/timecount_cnst[4] ), .S(\noisestate_0/N_228 ), 
        .Y(\noisestate_0/timecount_5[8] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[3] ));
    DFN1E1 \scalestate_0/timecount_ret_7  (.D(
        \scalestate_0/timecount_cnst_m_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_cnst_m_0_reto[3] ));
    DFN1E1 \top_code_0/noisedata[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[8] ));
    DFN1 \noisestate_0/CS[6]  (.D(\noisestate_0/CS_RNO[6]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[6]_net_1 ));
    AOI1D \timer_top_0/state_switch_0/dataout_RNO_5[6]  (.A(
        \scalestate_0/timecount_cnst_m_reto[6] ), .B(
        \scalestate_0/timecount_20_iv_10_reto[6] ), .C(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_213 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[3]  (.A(
        \timer_top_0/state_switch_0/N_227 ), .B(
        \timer_top_0/state_switch_0/N_229 ), .C(
        \timer_top_0/state_switch_0/N_228 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[3] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m134  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_131 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_134 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_135 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_62_i ));
    OR2 \scalestate_0/CS_RNIK8HJ[3]  (.A(\scalestate_0/CS[3]_net_1 ), 
        .B(\scalestate_0/CS[9]_net_1 ), .Y(\scalestate_0/N_1197 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI4AKD[1]  (.A(
        \sd_acq_top_0/count_10[1] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[1]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_6[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m278  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_275 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_278 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_279 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m140  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_139 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_140 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_141 ));
    AO1A \scalestate_0/timecount_ret_1_RNO_5  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[5]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[5] ), .Y(
        \scalestate_0/timecount_20_iv_1[5] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[14]  (.A(
        \scalestate_0_timecount[14] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_263 ));
    DFN1E1 \scalestate_0/timecount_ret_88  (.D(
        \scalestate_0/timecount_20_iv_6[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[10] ));
    MX2 \state_1ms_0/timecount_RNO_0[8]  (.A(
        \state_1ms_0/timecount_8[8] ), .B(\state_1ms_0_timecount[8] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_75 ));
    DFN1 \CAL_0/cal_div_0/count[5]  (.D(\CAL_0/cal_div_0/count_5[5] ), 
        .CLK(ddsclkout_c), .Q(\CAL_0/cal_div_0/count[5]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m157  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_154 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_157 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_158 ));
    XOR2 \PLUSE_0/qq_coder_1/un1_qq_para2_2[0]  (.A(
        \PLUSE_0/qq_para2[2] ), .B(\PLUSE_0/count_7[2] ), .Y(
        \PLUSE_0/qq_coder_1/un1_qq_para2_2[0]_net_1 ));
    OA1C \top_code_0/cal_load_RNO  (.A(\top_code_0/N_204 ), .B(
        top_code_0_cal_load), .C(\top_code_0/N_272 ), .Y(
        \top_code_0/N_64 ));
    MX2A \scalestate_0/reset_out_RNO_0  (.A(\scalestate_0/N_1097 ), .B(
        net_45), .S(\scalestate_0/N_1189 ), .Y(\scalestate_0/N_540 ));
    DFN1E1 \noisestate_0/dectime[10]  (.D(\top_code_0_noisedata[10] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \noisestate_0/dectime[10]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_128  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_128_Y ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/ADD_20x20_slow_I19_Y_0 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[19] ));
    NOR2B \pd_pluse_top_0/pd_pluse_coder_0/i_RNO[5]  (.A(net_27), .B(
        bri_dump_sw_0_tetw_pluse), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_0[5] ));
    NOR3B \DUMP_OFF_1/off_on_state_0/cs_RNO[1]  (.A(
        nsctrl_choice_0_dumponoff_rst), .B(\DUMP_OFF_1/i_4[0] ), .C(
        \DUMP_OFF_1/off_on_state_0/N_10 ), .Y(
        \DUMP_OFF_1/off_on_state_0/cs_nsss[1] ));
    OA1 \syn_md_module_1/syn_md_0/count_RNO_2[2]  (.A(
        \syn_md_module_1/syn_md_0/count[0]_net_1 ), .B(
        \syn_md_module_1/syn_md_0/count[1]_net_1 ), .C(
        \syn_md_module_1/syn_md_0/count[2]_net_1 ), .Y(
        \syn_md_module_1/syn_md_0/count_n2_i_a2_0 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i12_mux ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[16]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m43_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[16] ));
    DFN1E1 \top_code_0/dumpdata[4]  (.D(\GPMI_0_dataout_0[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[4] ));
    OR2B \DUMP_0/dump_state_0/cs_RNO_3[5]  (.A(
        \DUMP_0/dump_state_0/cs[4]_net_1 ), .B(\DUMP_0/i_0[3] ), .Y(
        \DUMP_0/dump_state_0/N_1497_tz_tz ));
    NOR3 \DDS_0/dds_state_0/para_RNO[18]  (.A(
        \DDS_0/dds_state_0/N_504 ), .B(\DDS_0/dds_state_0/N_503 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[18] ), .Y(
        \DDS_0/dds_state_0/N_163 ));
    DFN1E1 \top_code_0/plusedata[12]  (.D(\GPMI_0_dataout[12] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[12] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[21]  (.D(
        \top_code_0_dds_configdata[4] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[21]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m33  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_30 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_33 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_34 ));
    DFN1 \DDS_0/dds_state_0/cs[5]  (.D(
        \DDS_0/dds_state_0/cs_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[5]_net_1 ));
    AO1 \scalestate_0/timecount_ret_62_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[12]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[12] ), .Y(
        \scalestate_0/timecount_20_iv_4[12] ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_10  (.A(\xd_in[4] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[4] ));
    DFN1E1 \scanstate_0/dectime[11]  (.D(\top_code_0_scandata[11] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_0_sqmuxa_net_1 ), .Q(
        \scanstate_0/dectime[11]_net_1 ));
    OA1C \top_code_0/dumpload_RNO  (.A(\top_code_0/N_218 ), .B(
        top_code_0_dumpload), .C(\top_code_0/N_278 ), .Y(
        \top_code_0/N_70 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_11  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_93_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_41_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_11_Y ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_12_inst  (.A(
        \sd_acq_top_0/count_1[9] ), .B(\sd_acq_top_0/count_1[10] ), .C(
        \sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ));
    DFI0 \DSTimer_0/DFI0_1  (.D(\DSTimer_0/net_0 ), .CLK(GLA_net_1), 
        .QN(\DSTimer_0/DFI0_1_QN ));
    DFN1E1 \top_code_0/sigtimedata[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[15] ));
    DFN1 \state_1ms_0/timecount[9]  (.D(
        \state_1ms_0/timecount_RNO[9]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[9] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m53  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[9] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i16_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_54_i ));
    RAM512X18 #( .MEMORYFILE("RAM_R10C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R10C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_10_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_10_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_0_net )
        );
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[1]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n1 ));
    RAM512X18 #( .MEMORYFILE("RAM_R11C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R11C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_11_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_11_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_0_net )
        );
    MX2 \scanstate_0/timecount_1_RNO_0[3]  (.A(
        \scanstate_0/dectime[3]_net_1 ), .B(
        \scanstate_0/acqtime[3]_net_1 ), .S(\scanstate_0/CS[4]_net_1 ), 
        .Y(\scanstate_0/N_61 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[4]  (.D(
        \top_code_0_pd_pluse_data[4] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[4]_net_1 ));
    IOPAD_IN \xa_pad[3]/U0/U0  (.PAD(xa[3]), .Y(\xa_pad[3]/U0/NET1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m271  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_268 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_271 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_272 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI0E6C3[12]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_7[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_6[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_15[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_18[0] ));
    NOR3 \top_code_0/nstateload_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_160 ), .Y(
        \top_code_0/N_288 ));
    NOR3B \sd_acq_top_0/sd_sacq_timer_0/count_RNO[0]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/count_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[0] ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_0[0]  (.A(
        \sd_acq_top_0/count[21] ), .B(\sd_acq_top_0/count[17] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_0[0]_net_1 ));
    IOIN_IB \gpio_pad/U0/U1  (.YIN(\gpio_pad/U0/NET1 ), .Y(gpio_c));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/SAND2_27_inst  (
        .A(\sd_acq_top_0/count[18] ), .B(\sd_acq_top_0/count[19] ), .C(
        \sd_acq_top_0/count[20] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_33_net ));
    NOR3C 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa_0_a2  
        (.A(\top_code_0_pd_pluse_choice[0] ), .B(
        \top_code_0_pd_pluse_choice[1] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/N_12 ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/UXOR2_12_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_15_net ), 
        .B(\sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[15] ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[6]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[6] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count_3[6] ));
    XA1A \PLUSE_0/qq_coder_0/i_RNO_2[1]  (.A(\PLUSE_0/count_9[0] ), .B(
        \PLUSE_0/qq_para1[0] ), .C(\PLUSE_0/qq_coder_0/i_0_0[1] ), .Y(
        \PLUSE_0/qq_coder_0/i_0_2[1] ));
    IOPAD_TRI \sd_acq_en_pad/U0/U0  (.D(\sd_acq_en_pad/U0/NET1 ), .E(
        \sd_acq_en_pad/U0/NET2 ), .PAD(sd_acq_en));
    DFN1 \DUMP_0/dump_timer_0/count[7]  (.D(
        \DUMP_0/dump_timer_0/count_n7 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[7] ));
    DFN1 \DUMP_0/dump_timer_0/count[10]  (.D(
        \DUMP_0/dump_timer_0/count_n10 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count[10] ));
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/en_RNO  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0_en ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/en_RNO_0 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIE07K[7]  (.A(
        \sd_acq_top_0/count_3[7] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[7]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_5[0] ));
    DFN1E1 \scalestate_0/timecount_ret_48  (.D(
        \scalestate_0/timecount_20_0_iv_0[17] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_0_iv_0_reto[17] ));
    DFN1E1 \top_code_0/s_addchoice_3[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_3[4] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[3]  (.D(
        \top_code_0_state_1ms_data[3] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[3]_net_1 ));
    XOR2 \PLUSE_0/qq_coder_0/i_RNO_3[1]  (.A(\PLUSE_0/qq_para1[1] ), 
        .B(\PLUSE_0/count_9[1] ), .Y(
        \PLUSE_0/qq_coder_0/un1_count_1[0] ));
    NOR3 \pd_pluse_top_0/pd_pluse_state_0/en1_RNO_0  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_166 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_184 ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[7]  (.D(
        \DUMP_0/dump_coder_0/para5_4[7] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[7]_net_1 ));
    AX1C 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_ADD_20x20_slow_I19_Y  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[18] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_41_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[19] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/ADD_20x20_slow_I19_Y_3 )
        );
    DFN1E1 \scalestate_0/PLUSETIME90[9]  (.D(
        \top_code_0_scaledatain[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[9]_net_1 ));
    XO1 \scalestate_0/M_pulse_RNO_2  (.A(
        \scalestate_0/necount[4]_net_1 ), .B(
        \scalestate_0/M_NUM[4]_net_1 ), .C(\scalestate_0/M_pulse8_10 ), 
        .Y(\scalestate_0/M_pulse8_NE_4 ));
    IOPAD_IN \xa_pad[13]/U0/U0  (.PAD(xa[13]), .Y(\xa_pad[13]/U0/NET1 )
        );
    XOR2 \scalestate_0/M_pulse_RNO_11  (.A(
        \scalestate_0/M_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(\scalestate_0/M_pulse8_5 )
        );
    DFN1E1 \top_code_0/pd_pluse_choice[2]  (.D(\GPMI_0_dataout[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_choice_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_choice[2] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_RNO_net_1 )
        , .CLK(ddsclkout_c), .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/s_clk_div4_0/count_net_1 ));
    XA1 \DUMP_0/off_on_timer_1/count_RNO[2]  (.A(
        \DUMP_0/off_on_timer_1/count_c1 ), .B(\DUMP_0/count_0[2] ), .C(
        \DUMP_0/off_on_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/off_on_timer_1/count_n2 ));
    XA1 \DUMP_0/dump_timer_0/count_RNO[1]  (.A(\DUMP_0/count_1[1] ), 
        .B(\DUMP_0/count_1[0] ), .C(
        \DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_0/dump_timer_0/count_n1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[14]  (.D(
        \top_code_0_sd_sacq_data[14] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[14]_net_1 ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/en1  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/en1_RNO_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/en1_net_1 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[13]  (.D(
        \ClockManagement_0/long_timer_0/count_n13 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[13]_net_1 ));
    OR2B \DUMP_OFF_0/off_on_state_0/state_over_RNO  (.A(
        \DUMP_OFF_0/off_on_state_0/N_12_mux ), .B(
        bri_dump_sw_0_reset_out), .Y(\DUMP_OFF_0/off_on_state_0/N_9 ));
    NOR2A \scalestate_0/timecount_ret_58_RNO_2  (.A(
        \scalestate_0/S_DUMPTIME[0]_net_1 ), .B(\scalestate_0/N_1089 ), 
        .Y(\scalestate_0/S_DUMPTIME_m[0] ));
    AOI1D \scalestate_0/timecount_ret_4_RNO  (.A(\scalestate_0/N_1203 )
        , .B(\scalestate_0/CS[16]_net_1 ), .C(top_code_0_scale_rst_3), 
        .Y(\scalestate_0/timecount_cnst_m_0[2] ));
    NOR2B \DDS_0/dds_state_0/para_RNO_0[33]  (.A(
        \DDS_0/dds_state_0/para[34]_net_1 ), .B(
        \DDS_0/dds_state_0/N_534 ), .Y(\DDS_0/dds_state_0/N_522 ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNISPBI1[0]  (.A(
        \ClockManagement_0/clk_10k_0/count[7]_net_1 ), .B(
        \ClockManagement_0/clk_5M_en ), .C(
        \ClockManagement_0/clk_10k_0/count[0]_net_1 ), .Y(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_6 ));
    AO1B \PLUSE_0/qq_state_1/stateover_RNO  (.A(
        \PLUSE_0/qq_state_1_stateover ), .B(\PLUSE_0/qq_state_1/N_84 ), 
        .C(\PLUSE_0/qq_state_1/cs4 ), .Y(
        \PLUSE_0/qq_state_1/stateover_RNO_1 ));
    OA1B \PLUSE_0/bri_coder_0/bri_cycle  (.A(
        \PLUSE_0/bri_coder_0/un2lto7_2_net_1 ), .B(
        \PLUSE_0/bri_coder_0/un2lto7_3_net_1 ), .C(
        \PLUSE_0/bri_coder_0_half ), .Y(PLUSE_0_bri_cycle));
    AO1A \scalestate_0/timecount_ret_28_RNO_1  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[1]_net_1 ), 
        .C(\scalestate_0/PLUSETIME90_m[1] ), .Y(
        \scalestate_0/timecount_20_iv_1[1] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m212  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[9] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_213 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m71  (.A(
        \top_code_0_s_addchoice_0[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[6] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_72 ));
    NOR2B \plusestate_0/pluse_acq_RNO  (.A(\plusestate_0/N_122 ), .B(
        top_code_0_pluse_rst), .Y(\plusestate_0/pluse_acq_RNO_net_1 ));
    MX2B \top_code_0/dump_sustain_RNO_0  (.A(top_code_0_dump_sustain), 
        .B(\xa_c[0] ), .S(\top_code_0/N_262 ), .Y(\top_code_0/N_808 ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[10]  (.D(
        \top_code_0_state_1ms_data[10] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[10]_net_1 ));
    NOR3C \scalestate_0/un1_PLUSETIME9032_5_i_a2_0  (.A(
        top_code_0_scaleload), .B(\top_code_0_scalechoice_0[4] ), .C(
        \top_code_0_scalechoice_0[1] ), .Y(
        \scalestate_0/un1_PLUSETIME9032_5_i_a2_0_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[2]  (.D(\GPMI_0_dataout_0[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[2] ));
    NOR3 \top_code_0/scanload_RNO_1  (.A(\top_code_0/N_151 ), .B(
        \top_code_0/N_142 ), .C(\top_code_0/N_159 ), .Y(
        \top_code_0/N_308 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[7]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_58_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[7] ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[5]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c4 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n5 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[4]  (.D(
        \top_code_0_scaledatain[4] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[4]_net_1 ));
    DFN1 \top_code_0/state_1ms_rst_n_0_0  (.D(
        \top_code_0/state_1ms_rst_n_0_0_RNI848T5_net_1 ), .CLK(
        GLA_net_1), .Q(top_code_0_state_1ms_rst_n_0));
    DFN1E1 \top_code_0/cal_data[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[2] ));
    NOR2A \scalestate_0/timecount_RNO_4[21]  (.A(
        \scalestate_0/CUTTIME90[21]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[21] ));
    DFN1E0 \DDS_0/dds_state_0/para[9]  (.D(\DDS_0/dds_state_0/N_14 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[9]_net_1 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m36  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[13] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i22_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_37_i ));
    DFN1E1 \scalestate_0/PLUSETIME90[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[5]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_4  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR0_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR1_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_4_Y ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[4]  (.D(
        \top_code_0_bri_datain[14] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para3[4] ));
    DFN1 \timer_top_0/timer_0/timedata[0]  (.D(
        \timer_top_0/timer_0/timedata_4[0] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[0]_net_1 ));
    OR2A \DDS_0/dds_state_0/cs_RNO_0[1]  (.A(
        \DDS_0/dds_state_0/cs[1]_net_1 ), .B(\DDS_0/i[1] ), .Y(
        \DDS_0/dds_state_0/N_229 ));
    DFN1E1 \top_code_0/n_divnum[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[1] ));
    DFN1E1 \top_code_0/bri_datain[12]  (.D(\GPMI_0_dataout[12] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[12] ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNI4P6F3[11]  
        (.A(\pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_1[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_0[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_9[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_12[0] ));
    AO1C \plusestate_0/CS_RNO_0[2]  (.A(\plusestate_0/CS[1]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_srsts_i_0[2] ));
    NOR3C \scalestate_0/timecount_ret_59_RNO_3  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[0]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[0] ));
    NOR2B \scalestate_0/timecount_ret_46_RNO  (.A(
        \scalestate_0/OPENTIME_TEL[16]_net_1 ), .B(
        \scalestate_0/N_258_0 ), .Y(\scalestate_0/OPENTIME_TEL_m[16] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_58_i ));
    AND2 \bridge_div_0/dataall_1_I_6  (.A(\top_code_0_scaleddsdiv[2] ), 
        .B(\top_code_0_scaleddsdiv[5] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_g_array_0_2[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_40  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_20_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_52_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_40_Y ));
    DFN1 \DDS_0/dds_state_0/cs[2]  (.D(\DDS_0/dds_state_0/N_38 ), .CLK(
        GLA_net_1), .Q(\DDS_0/dds_state_0/cs[2]_net_1 ));
    RAM512X18 #( .MEMORYFILE("RAM_R14C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R14C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_14_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_14_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_10_net )
        , .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_9_net )
        , .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_8_net )
        , .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_7_net )
        , .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_6_net )
        , .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_5_net )
        , .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_4_net )
        , .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_3_net )
        , .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_2_net )
        , .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_1_net )
        , .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_0_net )
        );
    DFN1 \scalestate_0/strippluse[5]  (.D(
        \scalestate_0/strippluse_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[5] ));
    DFN1C0 \PLUSE_0/bri_coder_0/i[2]/U1  (.D(
        \PLUSE_0/bri_coder_0/i[2]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/i_3[2] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m154  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_155 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[17]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[17]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_498 ));
    DFN1E1 \scalestate_0/PLUSETIME90[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[11]_net_1 ));
    XOR2 \bridge_div_0/dataall_1_I_8  (.A(\top_code_0_scaleddsdiv[2] ), 
        .B(\top_code_0_scaleddsdiv[5] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_pog_array_0_1[0] ));
    DFN1 \PLUSE_0/qq_timer_1/count[3]  (.D(
        \PLUSE_0/qq_timer_1/count_n3 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_7[3] ));
    DFN1 \topctrlchange_0/soft_dump  (.D(
        \topctrlchange_0/soft_dump_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        soft_dump_net_0));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[9]  (
        .D(\s_acq_change_0_s_acqnum[9] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[9]_net_1 )
        );
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNIURCQ1[12]  (.A(
        \sd_acq_top_0/count_0[12] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[12]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_NE_7[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_165  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_148_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_6_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_165_Y ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[8]  (.D(
        \ClockManagement_0/long_timer_0/count_n8 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[8]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i22_mux ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNI8J6B[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[6]_net_1 ), .B(
        \sd_acq_top_0/count_3[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_6[0] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_8  (.A(
        \timer_top_0/dataout[14] ), .B(
        \timer_top_0/timer_0/timedata[14]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_8_Y ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m121  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[3] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_122 ));
    RAM512X18 #( .MEMORYFILE("RAM_R3C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R3C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_3_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_3_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_0_net ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_1_0_0_ADD_12x12_slow_I6_un1_CO1  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N152 ), 
        .B(\s_acq_change_0_s_stripnum[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I6_un1_CO1 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[7]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n7 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIS70P[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[10]_net_1 ), .B(
        \sd_acq_top_0/count_1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_10[0] ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[10]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[10] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[10] ));
    DFN1 \s_acq_change_0/s_acqnum[6]  (.D(
        \s_acq_change_0/s_acqnum_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[6] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_4  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m39 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[3] )
        );
    DFN1 \DDS_0/dds_timer_0/count[2]  (.D(\DDS_0/dds_timer_0/count_n2 )
        , .CLK(GLA_net_1), .Q(\DDS_0/count[2] ));
    NOR2B \DDS_0/dds_state_0/para_RNO_3[7]  (.A(
        \top_code_0_dds_configdata[6] ), .B(\DDS_0/dds_state_0/N_538 ), 
        .Y(\DDS_0/dds_state_0/N_270 ));
    NOR2 \DUMP_OFF_1/off_on_coder_0/i_RNO_0[1]  (.A(
        \DUMP_OFF_1/count_4[1] ), .B(\DUMP_OFF_1/count_4[0] ), .Y(
        \DUMP_OFF_1/off_on_coder_0/i_0_1[1] ));
    DFN1E0 \DUMP_0/dump_coder_0/para4[8]  (.D(
        \DUMP_0/dump_coder_0/para4_4[8]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_3_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para4[8]_net_1 ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_29  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m39 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[5] )
        );
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_38_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m44_5 ));
    NOR3B 
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa_0_a2  
        (.A(\top_code_0_pd_pluse_choice[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/N_12 ), .C(
        \top_code_0_pd_pluse_choice[1] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ));
    OA1A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[9]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs[9]_net_1 ), .B(
        \pd_pluse_top_0/i_1[2] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_i[0]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_177 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[11]  
        (.D(\s_acq_change_0_s_acqnum[11] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[11]_net_1 )
        );
    NOR2B \scalestate_0/necount_RNO[6]  (.A(\scalestate_0/N_736 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[6]_net_1 ));
    DFN1E1 \top_code_0/scandata[11]  (.D(\GPMI_0_dataout[11] ), .CLK(
        GLA_net_1), .E(\top_code_0/scandata_1_sqmuxa ), .Q(
        \top_code_0_scandata[11] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_137  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_137_Y ));
    DFN1E1 \scalestate_0/timecount_ret_68  (.D(
        \scalestate_0/timecount_20_iv_8[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[14] ));
    AND3 \scalestate_0/necount_inc_0/AND2_1_8_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount_inc_0/inc_5_net ), .C(
        \scalestate_0/necount_inc_0/inc_8_net ), .Y(
        \scalestate_0/necount_inc_0/Rcout_8_net ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m35  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_20 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_35 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_t[1] ));
    DFN1E1 \scalestate_0/CUTTIME90[18]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1701 ), .Q(\scalestate_0/CUTTIME90[18]_net_1 ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_4  (.A(
        \timer_top_0/timer_0/timedata[2]_net_1 ), .B(
        \timer_top_0/dataout[2] ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_4_Y ));
    IOTRI_OR_EB \Q1Q8_pad/U0/U1  (.D(
        \PLUSE_0/qq_state_0/Q1Q8_Q2Q7_RNO_net_1 ), .E(VCC), .OCLK(
        GLA_net_1), .DOUT(\Q1Q8_pad/U0/NET1 ), .EOUT(
        \Q1Q8_pad/U0/NET2 ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[5]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_14_1 ), .Y(
        \timer_top_0/timer_0/timedata_4[5] ));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_10  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[6] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_COMP0_E[1] )
        );
    CLKINT 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enadd_RNIH9JE_0  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/clk_add_i ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ));
    XOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNIAQ6E[2]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_12 ), 
        .B(\s_acq_change_0_s_stripnum[2] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[2]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_2 ));
    OR3 \scalestate_0/timecount_ret_57_RNO  (.A(
        \scalestate_0/CUTTIME180_m[0] ), .B(
        \scalestate_0/OPENTIME_m[0] ), .C(
        \scalestate_0/timecount_20_iv_3[0] ), .Y(
        \scalestate_0/timecount_20_iv_7[0] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_54  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_54_Y ));
    NOR2B \DDS_0/dds_state_0/para_reg_100_e_0  (.A(
        top_code_0_dds_choice), .B(top_code_0_dds_load), .Y(
        \DDS_0/dds_state_0/N_569_0 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m47  
        (.A(\s_acq_change_0_s_stripnum[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[8]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i14_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_48_i ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[1]  (
        .D(\top_code_0_s_periodnum[1] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[1]_net_1 )
        );
    DFN1 \scanstate_0/CS[4]  (.D(\scanstate_0/CS_RNO_2[4] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[4]_net_1 ));
    DFN1 \PLUSE_0/qq_timer_0/count[3]  (.D(
        \PLUSE_0/qq_timer_0/count_n3 ), .CLK(GLA_net_1), .Q(
        \PLUSE_0/count_9[3] ));
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[2]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[2]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 )
        );
    NOR2A \DUMP_0/dump_coder_0/para2_4[11]  (.A(
        \top_code_0_dumpdata_0[11] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[11]_net_1 ));
    XNOR2 \scalestate_0/necount_cmp_1/XNOR2_3  (.A(
        \scalestate_0/necount[8]_net_1 ), .B(
        \scalestate_0/NE_NUM[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/XNOR2_3_Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m308  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_305 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_308 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_309 ));
    AO1B \scalestate_0/CS_RNI44CR[20]  (.A(\scalestate_0/CS[20]_net_1 )
        , .B(top_code_0_scale_rst_1), .C(\scalestate_0/N_1093 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_6_0 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI9AN5[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_9[0] ));
    OA1C \top_code_0/acqclken_RNO  (.A(\top_code_0/N_199 ), .B(
        top_code_0_acqclken), .C(\top_code_0/N_268 ), .Y(
        \top_code_0/N_60 ));
    DFN1 \ClockManagement_0/clk_div500_0/count[0]  (.D(
        \ClockManagement_0/clk_div500_0/count_5[0] ), .CLK(GLA_net_1), 
        .Q(\ClockManagement_0/clk_div500_0/count[0]_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_4[11]  (.A(
        \state_1ms_0/S_DUMPTIME[11]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[11] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[11] ));
    IOBI_IB_OB_EB \xd_pad[7]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[7] ), .E(\GPMI_0.tri_state_0.xd_1 )
        , .YIN(\xd_pad[7]/U0/NET3 ), .DOUT(\xd_pad[7]/U0/NET1 ), .EOUT(
        \xd_pad[7]/U0/NET2 ), .Y(\xd_in[7] ));
    AO1 \scanstate_0/dumpoff_ctr_RNO_0  (.A(scanstate_0_dumpoff_ctr), 
        .B(\scanstate_0/N_255 ), .C(\scanstate_0/CS[5]_net_1 ), .Y(
        \scanstate_0/N_113 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m248  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_245 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_248 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_249 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m55  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[8] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i14_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_56_i ));
    NOR3C \scalestate_0/timecount_ret_60_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[12]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[12] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_120  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_8_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_8_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_120_Y ));
    XO1 \DUMP_0/dump_coder_0/para4_RNIK3651[9]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_coder_0/para4[9]_net_1 ), .C(
        \DUMP_0/dump_coder_0/un1_count_1_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_5[0] ));
    XO1 \DUMP_0/dump_coder_0/para4_RNI8N551[6]  (.A(
        \DUMP_0/count_0[6] ), .B(\DUMP_0/dump_coder_0/para4[6]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_1_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_1_NE_1[0] ));
    AO1 \state_1ms_0/timecount_RNO_2[0]  (.A(
        \state_1ms_0/M_DUMPTIME[0]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[0] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[0] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[7] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_58_i ));
    DFN1P0 \PLUSE_0/bri_state_0/cs[13]  (.D(
        \PLUSE_0/bri_state_0/cs_RNO[13]_net_1 ), .CLK(ddsclkout_c), 
        .PRE(\PLUSE_0/bri_state_0/en_net_1 ), .Q(
        \PLUSE_0/bri_state_0/cs_i_0[13] ));
    DFN1 \timer_top_0/timer_0/timedata[5]  (.D(
        \timer_top_0/timer_0/timedata_4[5] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[5]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[21]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_426 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[21]_net_1 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[8]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[8] ));
    DFN1E1 \top_code_0/scaledatain[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[2] ));
    NOR2B \topctrlchange_0/soft_dump_RNO  (.A(\topctrlchange_0/N_11 ), 
        .B(net_27), .Y(\topctrlchange_0/soft_dump_RNO_0_net_1 ));
    DFN1E1 \plusestate_0/DUMPTIME[8]  (.D(\top_code_0_plusedata[8] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[8]_net_1 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[6]  (.A(\DDS_0/dds_state_0/N_277 )
        , .B(\DDS_0/dds_state_0/N_276 ), .C(
        \DDS_0/dds_state_0/para_9_i_0_1[6] ), .Y(
        \DDS_0/dds_state_0/N_44 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[7]  (.D(
        \top_code_0_pd_pluse_data[7] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[7]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_2_RNO_3  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[6]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[6] ));
    OR2B \DUMP_ON_0/off_on_state_0/state_over_RNO  (.A(
        \DUMP_ON_0/off_on_state_0/N_12_mux ), .B(OR2_2_Y), .Y(
        \DUMP_ON_0/off_on_state_0/N_9 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[8]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[8] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[8] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[11]  (.A(
        \timer_top_0/state_switch_0/N_197 ), .B(
        \timer_top_0/state_switch_0/N_199 ), .C(
        \timer_top_0/state_switch_0/N_198 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[11] ));
    AO1C \plusestate_0/CS_RNO_0[5]  (.A(\plusestate_0/CS[9]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_srsts_i_0[5] ));
    NOR3C \ClockManagement_0/clk_10k_0/count_RNIMH9O1[3]  (.A(
        \ClockManagement_0/clk_10k_0/count[4]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/count[3]_net_1 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_2 ), .Y(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_5 ));
    IOPAD_IN \xa_pad[16]/U0/U0  (.PAD(xa[16]), .Y(\xa_pad[16]/U0/NET1 )
        );
    NOR2B \scalestate_0/timecount_ret_14_RNO_0  (.A(
        \scalestate_0/CUTTIME180_TEL[9]_net_1 ), .B(
        \scalestate_0/N_261 ), .Y(\scalestate_0/CUTTIME180_TEL_m[9] ));
    DFN1E1 \scalestate_0/OPENTIME[16]  (.D(\top_code_0_scaledatain[0] )
        , .CLK(GLA_net_1), .E(\scalestate_0/N_1681 ), .Q(
        \scalestate_0/OPENTIME[16]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNO[11]  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c10 ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n11 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNICJ09[9]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[9]_net_1 ), .B(
        \sd_acq_top_0/count_1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_9[0] ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[8]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[8] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_2_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ));
    NOR2A \scalestate_0/strippluse_RNO_1[4]  (.A(\scalestate_0/N_424 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(
        \scalestate_0/strippluse_6[4] ));
    AOI1B \DDS_0/dds_state_0/cs_RNO[1]  (.A(
        \DDS_0/dds_state_0/cs_i[0]_net_1 ), .B(
        \DDS_0/dds_state_0/N_229 ), .C(\DDS_0/dds_state_0/N_223 ), .Y(
        \DDS_0/dds_state_0/cs_RNO[1]_net_1 ));
    MX2 \s_acq_change_0/s_rst_RNO_0  (.A(\s_acq_change_0/s_rst_5 ), .B(
        s_acq_change_0_s_rst), .S(\top_code_0_change_0[1] ), .Y(
        \s_acq_change_0/N_68 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[0]_net_1 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_3  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[11]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_42_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[2] )
        );
    MX2 \state_1ms_0/timecount_RNO_0[10]  (.A(
        \state_1ms_0/timecount_8[10] ), .B(\state_1ms_0_timecount[10] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_77 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[3]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[3] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIA43I1[21]  (.A(
        \sd_acq_top_0/count[21] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[21]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_17[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_0[0] ));
    IOPAD_TRI \relay_on_pad[9]/U0/U0  (.D(\relay_on_pad[9]/U0/NET1 ), 
        .E(\relay_on_pad[9]/U0/NET2 ), .PAD(relay_on[9]));
    DFN1C0 \bridge_div_0/count[3]  (.D(\bridge_div_0/count_5[3] ), 
        .CLK(ddsclkout_c), .CLR(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[3]_net_1 ));
    MX2 \s_acq_change_0/s_stripnum_RNO_0[0]  (.A(
        \s_acq_change_0/s_stripnum_5[0] ), .B(
        \s_acq_change_0_s_stripnum[0] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_56 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m241  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_238 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_241 ), .S(
        \top_code_0_s_addchoice[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_242 ));
    OAI1 \scalestate_0/fst_lst_pulse_RNI3SS42  (.A(
        \scalestate_0/N_1209 ), .B(\scalestate_0/fst_lst_pulse_net_1 ), 
        .C(\scalestate_0/N_1196 ), .Y(\scalestate_0/un1_CS6_26_0 ));
    NOR2B \DDS_0/dds_timer_0/count_RNO[6]  (.A(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .B(
        \DDS_0/dds_timer_0/count_n6_tz ), .Y(
        \DDS_0/dds_timer_0/count_n6 ));
    DFN1E1 \scalestate_0/CUTTIME90[0]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[0]_net_1 ));
    DFN1E1 \scalestate_0/ACQ90_NUM[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ90_NUM[10]_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[7]  (
        .D(\s_acq_change_0_s_acqnum[7] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[7]_net_1 )
        );
    DFN1E1 \noisestate_0/acqtime[7]  (.D(\top_code_0_noisedata[7] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[7]_net_1 ));
    OA1B \top_code_0/pluse_lc_RNO  (.A(\top_code_0/N_160 ), .B(
        \top_code_0/N_175 ), .C(\top_code_0/N_291 ), .Y(
        \top_code_0/N_84 ));
    IOIN_IB \xa_pad[6]/U0/U1  (.YIN(\xa_pad[6]/U0/NET1 ), .Y(\xa_c[6] )
        );
    DFN1E1 \top_code_0/plusedata[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[8] ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_88_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/N_24 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 )
        , .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ));
    IOIN_IB \ADC_pad[10]/U0/U1  (.YIN(\ADC_pad[10]/U0/NET1 ), .Y(
        \ADC_c[10] ));
    IOTRI_OB_EB \relay_on_pad[7]/U0/U1  (.D(\relay_on_c[7] ), .E(VCC), 
        .DOUT(\relay_on_pad[7]/U0/NET1 ), .EOUT(
        \relay_on_pad[7]/U0/NET2 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[11]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[12]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_328 ));
    DFN1 \scalestate_0/pn_out  (.D(\scalestate_0/pn_out_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(scalestate_0_pn_out));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_2_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_2_net ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[0]  (.A(
        \timer_top_0/state_switch_0/N_240 ), .B(
        \timer_top_0/state_switch_0/N_241 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[0] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[0]_net_1 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m37  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_37_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[14]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/m37 ));
    MX2 \state1ms_choice_0/pluse_start_RNO_0  (.A(
        bri_dump_sw_0_off_test), .B(state_1ms_0_pluse_start), .S(
        top_code_0_state_1ms_start), .Y(
        \state1ms_choice_0/pluse_start_5 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[32]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[32]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_312 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[11]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[11] ));
    DFN1 \nsctrl_choice_0/sw_acq2  (.D(
        \nsctrl_choice_0/sw_acq2_RNO_0_net_1 ), .CLK(GLA_net_1), .Q(
        nsctrl_choice_0_sw_acq2));
    NOR2A \DUMP_0/dump_coder_0/para4_4[7]  (.A(
        \top_code_0_dumpdata_0[7] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[7]_net_1 ));
    AO1 \scalestate_0/timecount_ret_29_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[1]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[1] ), .Y(
        \scalestate_0/timecount_20_iv_4[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m7  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_6_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_7_0 ), .S(
        \top_code_0_s_addchoice_1[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_8_0 ));
    DFN1 \s_acq_change_0/s_stripnum[6]  (.D(
        \s_acq_change_0/s_stripnum_RNO[6]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[6] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/HND2_13_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_17_net ), .B(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_16_net ), .C(
        \sd_acq_top_0/count_0[12] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_13_net ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNIGT6S[2]  (
        .A(\pd_pluse_top_0/count_6[2] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[2]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_12[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_NE_4[0] ));
    XA1A \DSTimer_0/dump_sustain_timer_0/start_RNO_0  (.A(
        \DSTimer_0/dump_sustain_timer_0/count[3]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/data[3]_net_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/enable_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/start11_0 ));
    DFN1E1 \top_code_0/s_acqnum[8]  (.D(\GPMI_0_dataout[8] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[8] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_24  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR12_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR13_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_24_Y ));
    DFN1E0 \DDS_0/dds_state_0/para[3]  (.D(\DDS_0/dds_state_0/N_157 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[3]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI78N5[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[8]_net_1 ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_8[0] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m129  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[3] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_130 ));
    AO1C \scalestate_0/necount_cmp_1/AO1C_2  (.A(
        \scalestate_0/necount[4]_net_1 ), .B(
        \scalestate_0/NE_NUM[4]_net_1 ), .C(
        \scalestate_0/necount[3]_net_1 ), .Y(
        \scalestate_0/necount_cmp_1/AO1C_2_Y ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[19]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[19]_net_1 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI56N5[7]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[7]_net_1 ), .B(
        \sd_acq_top_0/count_3[7] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_7[0] ));
    NOR2A \plusestate_0/timecount_1_RNO[10]  (.A(\plusestate_0/N_81 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[10] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[6] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_60_i ));
    MX2 \scalestate_0/necount_RNO_0[10]  (.A(
        \scalestate_0/necount1[10] ), .B(
        \scalestate_0/necount[10]_net_1 ), .S(\scalestate_0/N_1179 ), 
        .Y(\scalestate_0/N_740 ));
    NOR2B \state_1ms_0/timecount_RNO_5[4]  (.A(
        \state_1ms_0/PLUSECYCLE[4]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[4] ));
    MX2 \scalestate_0/sw_acq2_RNO_0  (.A(\scalestate_0/N_1251_1 ), .B(
        scalestate_0_sw_acq2), .S(\scalestate_0/un1_CS6_34 ), .Y(
        \scalestate_0/N_541 ));
    DFN1 \s_acq_change_0/s_rst  (.D(\s_acq_change_0/s_rst_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(\s_acq_change_0/s_rst_net_1 ));
    AOI1A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_32  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[3] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[4] ), 
        .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT3_E[5] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_CMPLE_PO2_DWACT_COMP0_E[0] )
        );
    MX2 \scalestate_0/necount_RNO_0[9]  (.A(\scalestate_0/necount1[9] )
        , .B(\scalestate_0/necount[9]_net_1 ), .S(
        \scalestate_0/N_1179 ), .Y(\scalestate_0/N_739 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[10]_net_1 ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[11]  (.A(
        \scalestate_0/s_acqnum_7[11] ), .B(\scalestate_0_s_acqnum[11] )
        , .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_558 ));
    NOR2B \scalestate_0/load_out_RNO  (.A(\scalestate_0/N_572 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/load_out_RNO_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[14]  (.D(
        \top_code_0_dds_configdata[13] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[14]_net_1 ));
    AND3 \bridge_div_0/count_5_I_8  (.A(
        \bridge_div_0/count_RNIEMOM7[0]_net_1 ), .B(
        \bridge_div_0/count_RNIFNOM7[1]_net_1 ), .C(
        \bridge_div_0/count_RNIGOOM7[2]_net_1 ), .Y(\bridge_div_0/N_4 )
        );
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/cs[3]  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[3]_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0/cs[3]_net_1 )
        );
    DFN1E1 \scalestate_0/CUTTIME180_Tini[19]  (.D(
        \top_code_0_scaledatain[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[19]_net_1 ));
    OR3 \state_1ms_0/timecount_RNO_1[4]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[4] ), .B(
        \state_1ms_0/CUTTIME_m[4] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[4] ), .Y(
        \state_1ms_0/timecount_8[4] ));
    NOR2B \scalestate_0/strippluse_RNO[6]  (.A(\scalestate_0/N_565 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[6]_net_1 ));
    IOTRI_OB_EB \relay_close_pad[3]/U0/U1  (.D(\relay_close_c[3] ), .E(
        VCC), .DOUT(\relay_close_pad[3]/U0/NET1 ), .EOUT(
        \relay_close_pad[3]/U0/NET2 ));
    DFN1E1 \scalestate_0/ACQ180_NUM[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQ180_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQ180_NUM[10]_net_1 ));
    OR2 \scalestate_0/CS_RNI75VB[17]  (.A(\scalestate_0/CS[7]_net_1 ), 
        .B(\scalestate_0/CS[17]_net_1 ), .Y(\scalestate_0/N_1194 ));
    IOTRI_OB_EB \relay_close_pad[4]/U0/U1  (.D(\relay_close_c[4] ), .E(
        VCC), .DOUT(\relay_close_pad[4]/U0/NET1 ), .EOUT(
        \relay_close_pad[4]/U0/NET2 ));
    XA1 \DUMP_ON_0/off_on_timer_0/count_RNO[2]  (.A(
        \DUMP_ON_0/off_on_timer_0/count_c1 ), .B(
        \DUMP_ON_0/count_5[2] ), .C(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_n2 ));
    MX2C \DUMP_ON_0/off_on_state_0/cs_RNO_0[1]  (.A(
        \DUMP_ON_0/off_on_state_0/cs[1]_net_1 ), .B(\DUMP_ON_0/i_5[1] )
        , .S(DUMP_ON_0_dump_on), .Y(\DUMP_ON_0/off_on_state_0/N_10 ));
    DFN1E1 \top_code_0/scaledatain_0[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain_0[2] ));
    OAI1 \state_1ms_0/CS_i_RNO_0[0]  (.A(timer_top_0_clk_en_st1ms), .B(
        \state_1ms_0/CS_i[0]_net_1 ), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/N_204s_i_i_0 ));
    DFN1E1 \plusestate_0/timecount_1[8]  (.D(
        \plusestate_0/timecount_5[8] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[8] ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[3]  (
        .D(\top_code_0_s_periodnum[3] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/datareg[3]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m41  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_40 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_41 ), .S(
        \top_code_0_s_addchoice_0[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_42 ));
    NOR3C \timer_top_0/timer_0/time_up_RNO  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/cmp_result ), .Y(
        \timer_top_0/timer_0/time_up_RNO_net_1 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[4]  (.D(
        \top_code_0_state_1ms_data[4] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[4]_net_1 ));
    DFN1E1 \state_1ms_0/CUTTIME[6]  (.D(\top_code_0_state_1ms_data[6] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[6]_net_1 ));
    AND2 \timer_top_0/timer_0/un2_timedata_I_15  (.A(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .B(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .Y(
        \timer_top_0/timer_0/DWACT_FINC_E[1] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[6]  (.A(
        \plusestate_0_timecount[6] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_214 ));
    NOR3A \top_code_0/scanchoice_RNO_1  (.A(\top_code_0/N_329 ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_142 ), .Y(
        \top_code_0/N_306 ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[5]  (.A(
        \timer_top_0/state_switch_0/N_215 ), .B(
        \timer_top_0/state_switch_0/N_216 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[5] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[5]_net_1 ));
    AO1C \plusestate_0/timecount_1_RNO_1[5]  (.A(
        \plusestate_0/CS[4]_net_1 ), .B(\plusestate_0/N_303 ), .C(
        top_code_0_pluse_rst_0), .Y(\plusestate_0/N_251 ));
    DFN1E0 \DDS_0/dds_state_0/para[0]  (.D(\DDS_0/dds_state_0/N_203 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[0]_net_1 ));
    NOR3B \top_code_0/scaleddsdiv_1_sqmuxa_0_a2  (.A(
        \top_code_0/N_331 ), .B(\top_code_0/N_334 ), .C(
        \top_code_0/N_157 ), .Y(\top_code_0/scaleddsdiv_1_sqmuxa ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_33  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR14_7_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR15_7_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_4_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_33_Y ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[19]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[19] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[19] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[6]  (.D(
        \top_code_0_halfdata_0[6] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[6] ));
    NOR2B \top_code_0/relay_close_RNO[6]  (.A(\top_code_0/N_825 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[6]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m172  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_169 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_172 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_173 ));
    AND2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y ));
    DFN1 \DUMP_0/dump_state_0/cs[1]  (.D(
        \DUMP_0/dump_state_0/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[1]_net_1 ));
    DFN1 \top_code_0/state_1ms_start_ret_1  (.D(net_27), .CLK(
        GLA_net_1), .Q(\top_code_0/net_27_reto ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[10]_net_1 ));
    DFN1C0 \bridge_div_0/count[5]  (.D(\bridge_div_0/count_5[5] ), 
        .CLK(ddsclkout_c), .CLR(bri_dump_sw_0_reset_out), .Q(
        \bridge_div_0/count[5]_net_1 ));
    MX2B \scanstate_0/timecount_1_RNO[3]  (.A(\scanstate_0/N_61 ), .B(
        \scanstate_0/N_196 ), .S(\scanstate_0/N_233 ), .Y(
        \scanstate_0/timecount_5[3] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_2_Y ));
    DFN1E1 \scalestate_0/ACQTIME[5]  (.D(\top_code_0_scaledatain[5] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[5]_net_1 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[27]  (.A(
        \DDS_0/dds_state_0/N_476 ), .B(\DDS_0/dds_state_0/N_475 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[27] ), .Y(
        \DDS_0/dds_state_0/N_127 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[23]  (.A(
        \DDS_0/dds_state_0/N_301 ), .B(\DDS_0/dds_state_0/N_300 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[23] ), .Y(
        \DDS_0/dds_state_0/N_20 ));
    DFN1E1 \state_1ms_0/PLUSETIME[3]  (.D(
        \top_code_0_state_1ms_data[3] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[3]_net_1 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m160  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[2] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_161 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI02EB[0]  (.A(
        \sd_acq_top_0/count_10[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[0]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_9[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_7[0] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[7]  (.A(
        \timer_top_0/state_switch_0/N_205 ), .B(
        \timer_top_0/state_switch_0/N_206 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[7] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[7]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[11]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_50_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[11] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[8]  (.A(\DDS_0/dds_state_0/N_285 )
        , .B(\DDS_0/dds_state_0/N_284 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[8] ), .Y(
        \DDS_0/dds_state_0/N_12 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/i_RNO_24[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[15]_net_1 ), .B(
        \sd_acq_top_0/count_0[15] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_15[0] ));
    AO1 \state_1ms_0/timecount_RNO_4[15]  (.A(
        \state_1ms_0/S_DUMPTIME[15]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[15] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[15] ));
    DFN1 \scanstate_0/CS[2]  (.D(\scanstate_0/CS_RNO_2[2] ), .CLK(
        GLA_net_1), .Q(\scanstate_0/CS[2]_net_1 ));
    NOR3A \scalestate_0/necount_cmp_0/NOR3A_2  (.A(
        \scalestate_0/necount_cmp_0/OR2A_1_Y ), .B(
        \scalestate_0/necount_cmp_0/AO1C_0_Y ), .C(
        \scalestate_0/M_NUM[0]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/NOR3A_2_Y ));
    XA1 \DUMP_OFF_0/off_on_timer_0/count_RNO[2]  (.A(
        \DUMP_OFF_0/off_on_timer_0/count_c1 ), .B(
        \DUMP_OFF_0/count_3[2] ), .C(
        \DUMP_OFF_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_OFF_0/off_on_timer_0/count_n2 ));
    NOR2B \scalestate_0/necount_RNO[1]  (.A(\scalestate_0/N_731 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[1]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_14_RNO_3  (.A(
        \scalestate_0/OPENTIME[9]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[9] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[7]  (.D(
        \top_code_0_dds_configdata[6] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[7]_net_1 ));
    AO1C \scanstate_0/CS_RNO_0[6]  (.A(\scanstate_0/CS[5]_net_1 ), .B(
        timer_top_0_clk_en_scan), .C(net_33), .Y(
        \scanstate_0/CS_srsts_i_0[6] ));
    DFN1E1 \scalestate_0/timecount_ret_29  (.D(
        \scalestate_0/timecount_20_iv_8[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[1] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[13]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[14]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_337 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[2]  (.A(\DDS_0/dds_state_0/N_488 )
        , .B(\DDS_0/dds_state_0/N_487 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[2] ), .Y(
        \DDS_0/dds_state_0/N_155 ));
    DFN1 \top_code_0/noise_start_ret_3  (.D(\top_code_0/N_114 ), .CLK(
        GLA_net_1), .Q(\top_code_0/N_114_reto ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[8]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[9]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_285 ));
    DFN1E1 \scalestate_0/CUTTIME90[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1685 ), .Q(\scalestate_0/CUTTIME90[3]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[11]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[11] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_50_i ));
    XOR2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNO[7]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c6 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n7 ));
    OR2 \sd_acq_top_0/sd_sacq_state_0/en2_RNIG9AD  (.A(
        \sd_acq_top_0/sd_sacq_state_0/en2_net_1 ), .B(
        \sd_acq_top_0/sd_sacq_state_0/en1 ), .Y(sd_acq_en_c));
    DFN1E1 \scalestate_0/timecount_ret_34  (.D(
        \scalestate_0/timecount_20_iv_6[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[9] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[10]  (.A(\scalestate_0/N_458 ), 
        .B(\scalestate_0/ACQECHO_NUM[10]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[10] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[0]  (.D(
        \top_code_0_bri_datain[10] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para3[0] ));
    AND2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[11] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[10]  (.A(\scalestate_0/N_557 ), 
        .B(top_code_0_scale_rst_4), .Y(
        \scalestate_0/s_acqnum_1_RNO[10]_net_1 ));
    NOR3C \ClockManagement_0/clk_10k_0/count_RNI8ESK4[0]  (.A(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_5 ), .B(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_4 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa_6 ), .Y(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ));
    MX2 \top_code_0/relay_close_RNO_0[6]  (.A(\relay_close_c[6] ), .B(
        \GPMI_0_dataout[6] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_825 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[4]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[4] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[4] ));
    NOR2A \DDS_0/dds_state_0/para_reg_69_e_0  (.A(top_code_0_dds_load), 
        .B(top_code_0_dds_choice), .Y(\DDS_0/dds_state_0/N_538_0 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[2]  (.D(
        \DUMP_0/dump_coder_0/para2_4[2]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[2]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_64_i ));
    DFN1E1 \top_code_0/s_periodnum[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_periodnum_1_sqmuxa ), .Q(
        \top_code_0_s_periodnum[0] ));
    NOR3A \ClockManagement_0/long_timer_0/timeup_RNO_2  (.A(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_6 ), .B(
        \ClockManagement_0/long_timer_0/clear_n4_8 ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_9 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_11 ));
    AO18 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m25  
        (.A(\s_acq_change_0_s_stripnum[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[8]_net_1 )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i16_mux )
        );
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafive[4]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_0_net_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[4] ));
    OR3 \scalestate_0/timecount_ret_29_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[1] ), .B(
        \scalestate_0/OPENTIME_TEL_m[1] ), .C(
        \scalestate_0/timecount_20_iv_4[1] ), .Y(
        \scalestate_0/timecount_20_iv_8[1] ));
    OA1 \PLUSE_0/bri_state_0/cs_RNIT2MF1[1]  (.A(
        \PLUSE_0/bri_state_0/cs[1]_net_1 ), .B(
        \PLUSE_0/bri_state_0/N_179 ), .C(\PLUSE_0/i_3[2] ), .Y(
        \PLUSE_0/bri_state_0/N_180 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[10]  (.A(
        \DDS_0/dds_state_0/N_293 ), .B(\DDS_0/dds_state_0/N_292 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[10] ), .Y(
        \DDS_0/dds_state_0/N_16 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[11]  (.D(
        \top_code_0_dds_configdata[10] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[11]_net_1 ));
    AO1A \scalestate_0/timecount_ret_40_RNO  (.A(\scalestate_0/N_1089 )
        , .B(\scalestate_0/S_DUMPTIME[2]_net_1 ), .C(
        \scalestate_0/timecount_20_iv_1[2] ), .Y(
        \scalestate_0/timecount_20_iv_6[2] ));
    IOIN_IB \xa_pad[3]/U0/U1  (.YIN(\xa_pad[3]/U0/NET1 ), .Y(\xa_c[3] )
        );
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i14_mux ));
    MX2C \scalestate_0/s_acq180_RNO_2  (.A(\scalestate_0/CS[10]_net_1 )
        , .B(\scalestate_0/fst_lst_pulse_net_1 ), .S(
        \scalestate_0/CS[9]_net_1 ), .Y(\scalestate_0/un1_CS6_0 ));
    MX2 \top_code_0/relay_close_RNO_0[2]  (.A(\relay_close_c[2] ), .B(
        \GPMI_0_dataout_0[2] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_821 ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datafour[6]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafive_2_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[6] ));
    NOR3C \scalestate_0/timecount_ret_82_RNO_0  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[4]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[4] ));
    DFN1E1 \top_code_0/dds_configdata[3]  (.D(\GPMI_0_dataout[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[3] ));
    NOR2B \state_1ms_0/timecount_RNO[10]  (.A(\state_1ms_0/N_77 ), .B(
        top_code_0_state_1ms_rst_n_0), .Y(
        \state_1ms_0/timecount_RNO[10]_net_1 ));
    DFN1 \dds_change_0/dds_conf  (.D(\dds_change_0/dds_conf_RNO_net_1 )
        , .CLK(GLA_net_1), .Q(dds_change_0_dds_conf));
    OR3 \timer_top_0/state_switch_0/state_start_RNO  (.A(
        \timer_top_0/state_switch_0/N_295 ), .B(
        \timer_top_0/state_switch_0/N_296 ), .C(
        \timer_top_0/state_switch_0/state_start5_0_0_1 ), .Y(
        \timer_top_0/state_switch_0/state_start5 ));
    DFN1E1 \plusestate_0/DUMPTIME[9]  (.D(\top_code_0_plusedata[9] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[9]_net_1 ));
    NOR2A \scalestate_0/timecount_ret_82_RNO_1  (.A(
        \scalestate_0/DUMPTIME[4]_net_1 ), .B(\scalestate_0/N_1093 ), 
        .Y(\scalestate_0/DUMPTIME_m[4] ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_5_Y ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIQ70I[3]  (.A(
        \sd_acq_top_0/count_10[3] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[3]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_0[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_10[0] ));
    OR2A \top_code_0/scan_rst_RNIMNCI3  (.A(net_27), .B(
        \top_code_0/N_803 ), .Y(\top_code_0/scan_rst_RNIMNCI3_net_1 ));
    NOR2B \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_RNO  
        (.A(XRD_c), .B(n_acq_change_0_n_rst_n), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/clk_reg1_RNO_net_1 )
        );
    NOR2B \state_1ms_0/timecount_RNO_1[16]  (.A(
        \state_1ms_0/CUTTIME[16]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 )
        , .Y(\state_1ms_0/timecount_8[16] ));
    OR2 \top_code_0/un1_state_1ms_rst_n117_43_i_o2_1  (.A(
        \top_code_0/N_150 ), .B(\xa_c[1] ), .Y(\top_code_0/N_190 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m47  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[12] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/m47_0 ));
    OR2B \scalestate_0/CS_RNIR4SG[12]  (.A(\scalestate_0/CS[12]_net_1 )
        , .B(scalestate_0_ne_le), .Y(\scalestate_0/N_1195 ));
    OR3 \scalestate_0/timecount_ret_41_RNO  (.A(
        \scalestate_0/timecount_20_iv_0[2] ), .B(
        \scalestate_0/OPENTIME_TEL_m[2] ), .C(
        \scalestate_0/timecount_20_iv_4[2] ), .Y(
        \scalestate_0/timecount_20_iv_8[2] ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[31]  (.D(
        \top_code_0_dds_configdata[14] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_569_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[31]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_20  (.A(
        \timer_top_0/timer_0/N_16 ), .B(
        \timer_top_0/timer_0/timedata[7]_net_1 ), .Y(
        \timer_top_0/timer_0/I_20_0 ));
    NOR2B \DDS_0/dds_state_0/N_409_i_i_o2  (.A(\DDS_0/i[0] ), .B(
        dds_change_0_dds_rst), .Y(\DDS_0/dds_state_0/N_223 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNICO0P[18]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[18]_net_1 ), .B(
        \sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_18[0] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_15_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_1_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_15_net ));
    XOR2 \scalestate_0/fst_lst_pulse_RNO_10  (.A(
        \scalestate_0/NE_NUM[1]_net_1 ), .B(
        \scalestate_0/necount[1]_net_1 ), .Y(
        \scalestate_0/fst_lst_pulse8_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datatwo[1]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datatwo ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[1] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO[3]  (.A(
        \timer_top_0/state_switch_0/N_225 ), .B(
        \timer_top_0/state_switch_0/N_226 ), .C(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[3] ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[3]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1729 ), .Q(
        \scalestate_0/CUTTIME180_Tini[1]_net_1 ));
    DFN1E1 \top_code_0/state_1ms_data[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[3] ));
    DFN1E1 \top_code_0/noisedata[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[1] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[13]_net_1 ));
    NOR3C \scalestate_0/timecount_ret_77_RNO_3  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[6]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[6] ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[7]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[7] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[7] ));
    XA1C \ClockManagement_0/long_timer_0/timeup_RNO_10  (.A(
        \ClockManagement_0/long_timer_0/count[12]_net_1 ), .B(
        \top_code_0_sigtimedata[12] ), .C(
        \ClockManagement_0/long_timer_0/clear_n4_14 ), .Y(
        \ClockManagement_0/long_timer_0/timeup_0_sqmuxa_2 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m196  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_193 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_196 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_197 ));
    OR3 \DUMP_0/dump_coder_0/para3_RNI08LG6[10]  (.A(
        \DUMP_0/dump_coder_0/un1_count_2_NE_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_2_NE_6[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE[0] ));
    NOR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIEICT9[2]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_NE ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_11 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[9]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[9] ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/YAND2BB_21_inst  
        (.A(\sd_acq_top_0/count_1[9] ), .B(\sd_acq_top_0/count_1[10] ), 
        .C(\sd_acq_top_0/count_1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_16_net ));
    NOR2B \scalestate_0/CS_RNO[1]  (.A(\scalestate_0/N_1217 ), .B(
        top_code_0_scale_rst_3), .Y(\scalestate_0/CS_RNO_1[1] ));
    NOR2B \PLUSE_0/qq_coder_1/i_RNO[0]  (.A(\PLUSE_0/down ), .B(
        bri_dump_sw_0_reset_out), .Y(\PLUSE_0/qq_coder_1/i_RNO_8[0] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_9  (.A(
        \timer_top_0/dataout[19] ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_9_Y ));
    MX2 \state_1ms_0/timecount_RNO_0[13]  (.A(
        \state_1ms_0/timecount_8[13] ), .B(\state_1ms_0_timecount[13] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_80 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_15  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_6_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_6_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_12_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_15_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_19  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR4_3_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR5_3_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_13_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_19_Y ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9]/U0  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9] ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_n9 ), 
        .S(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/I_45 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[9]/Y ));
    DFN1E1 \scalestate_0/timecount_ret_8  (.D(
        \scalestate_0/timecount_20_iv_7[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[3] ));
    DFN1E1 \noisestate_0/acqtime[8]  (.D(\top_code_0_noisedata[8] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[8]_net_1 ));
    NOR3 \state_1ms_0/soft_dump_RNO_1  (.A(\state_1ms_0/CS[8]_net_1 ), 
        .B(\state_1ms_0/CS[1]_net_1 ), .C(\state_1ms_0/CS[2]_net_1 ), 
        .Y(\state_1ms_0/N_255 ));
    NOR3A \DUMP_0/dump_state_0/cs_RNO_1[5]  (.A(
        \DUMP_0/dump_state_0/N_1497_tz_tz ), .B(
        \DUMP_0/dump_state_0_on_start ), .C(
        \DUMP_0/dump_state_0/cs[6]_net_1 ), .Y(
        \DUMP_0/dump_state_0/cs_RNO_1[5]_net_1 ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIHHP03[6]  (.A(
        \ClockManagement_0/long_timer_0/count_c5 ), .B(
        \ClockManagement_0/long_timer_0/count[6]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_c6 ));
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_11_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_14_net ), .B(
        \sd_acq_top_0/count_0[14] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[14] ));
    IOIN_IB \ADC_pad[7]/U0/U1  (.YIN(\ADC_pad[7]/U0/NET1 ), .Y(
        \ADC_c[7] ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[11]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[4] ));
    DFN1 \state_1ms_0/CS[7]  (.D(\state_1ms_0/CS_RNO_3[7] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[7]_net_1 ));
    DFN1E1 \top_code_0/plusedata[14]  (.D(\GPMI_0_dataout[14] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[14] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[1]  (.D(
        \top_code_0_state_1ms_data[1] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[1]_net_1 ));
    AX1A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m4  (.A(
        \top_code_0_s_addchoice_0[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_313 ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signal_data_en[0] ));
    NOR3 \DDS_0/dds_state_0/para_RNO[22]  (.A(
        \DDS_0/dds_state_0/N_269 ), .B(\DDS_0/dds_state_0/N_460 ), .C(
        \DDS_0/dds_state_0/para_9_i_0_1[22] ), .Y(
        \DDS_0/dds_state_0/N_40 ));
    DFN1 \state_1ms_0/CS[8]  (.D(\state_1ms_0/CS_RNO_1[8] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[8]_net_1 ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[10]  (.D(
        \top_code_0_scaledatain[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[10]_net_1 ));
    NOR3C \DUMP_0/dump_timer_0/count_0_sqmuxa  (.A(
        \DUMP_0/dump_state_0_timer_start ), .B(
        state1ms_choice_0_dump_start), .C(state1ms_choice_0_reset_out), 
        .Y(\DUMP_0/dump_timer_0/count_0_sqmuxa_net_1 ));
    DFN1E1 \top_code_0/scaledatain[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[4] ));
    NOR2A \scalestate_0/timecount_ret_35_RNO_1  (.A(
        \scalestate_0/CUTTIME90[9]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[9] ));
    AO1 \scalestate_0/timecount_ret_22_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL[10]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[10] )
        , .Y(\scalestate_0/timecount_20_iv_3[10] ));
    OR2 \top_code_0/s_load_RNO_0  (.A(\top_code_0/N_192 ), .B(
        \top_code_0/N_150 ), .Y(\top_code_0/N_196 ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNI8DFH[0]  (.A(
        \DUMP_0/dump_coder_0/para3[0]_net_1 ), .B(\DUMP_0/count_1[0] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_0_0[0] ));
    XOR2 \bridge_div_0/dataall_1_I_9  (.A(\top_code_0_scaleddsdiv[0] ), 
        .B(\top_code_0_scaleddsdiv[3] ), .Y(
        \bridge_div_0/DWACT_ADD_CI_0_partial_sum[0] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_6_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_7_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_6_net ));
    DFN1E1 \scalestate_0/timecount_ret_70  (.D(
        \scalestate_0/timecount_20_iv_6[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[15] ));
    MX2 \PLUSE_0/bri_state_0/cs_RNO[13]  (.A(
        \PLUSE_0/bri_state_0/cs_i_0[13] ), .B(
        \PLUSE_0/bri_state_0/cs_i_0[12] ), .S(clk_4f_en), .Y(
        \PLUSE_0/bri_state_0/cs_RNO[13]_net_1 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_11_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_5_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_11_net ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[15]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/i_RNO[8]  (.A(
        state1ms_choice_0_reset_out), .B(
        \DUMP_0/dump_coder_0/i_reg16_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO[8]_net_1 ));
    DFN1E1 \top_code_0/sd_sacq_data[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m210  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_209 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_210 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_211 ));
    NOR2A \scalestate_0/timecount_ret_50_RNO_3  (.A(
        \scalestate_0/CUTTIME90[17]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[17] ));
    AND2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2_14_inst  (.A(
        \sd_acq_top_0/count_0[12] ), .B(\sd_acq_top_0/count_0[13] ), 
        .Y(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_20_net ));
    IOTRI_OB_EB \relay_on_pad[4]/U0/U1  (.D(\relay_on_c[4] ), .E(VCC), 
        .DOUT(\relay_on_pad[4]/U0/NET1 ), .EOUT(
        \relay_on_pad[4]/U0/NET2 ));
    OR2B \plusestate_0/CS_RNIL3FD[5]  (.A(\plusestate_0/CS[5]_net_1 ), 
        .B(top_code_0_pluse_rst), .Y(\plusestate_0/N_213 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m28  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i16_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[9] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i18_mux ));
    DFN1 \DUMP_0/dump_coder_0/i[5]  (.D(
        \DUMP_0/dump_coder_0/i_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i[5] ));
    DFN1E1 \scalestate_0/timecount_ret_4  (.D(
        \scalestate_0/timecount_cnst_m_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_cnst_m_0_reto[2] ));
    IOTRI_OB_EB \relay_on_pad[3]/U0/U1  (.D(\relay_on_c[3] ), .E(VCC), 
        .DOUT(\relay_on_pad[3]/U0/NET1 ), .EOUT(
        \relay_on_pad[3]/U0/NET2 ));
    OR3 \dds_change_0/dds_conf_RNO_1  (.A(\dds_change_0/dds_confin2_m )
        , .B(\dds_change_0/dds_confin3_m ), .C(
        \dds_change_0/dds_confin1_m ), .Y(\dds_change_0/dds_conf_6 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[9]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[9] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[9] ));
    NOR2A \PLUSE_0/bri_coder_0/half_0_I_7  (.A(\PLUSE_0/count_2[5] ), 
        .B(\PLUSE_0/half_para[5] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[0] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_6[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_66_i ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m101  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[4] ), .C(
        \top_code_0_s_addchoice_0[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_102 ));
    DFN1 \scalestate_0/strippluse[11]  (.D(
        \scalestate_0/strippluse_RNO[11]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[11] ));
    NOR2B \timer_top_0/state_switch_0/clk_en_pluse_0_0_a6_0_a2  (.A(
        top_code_0_pluse_str), .B(net_27), .Y(
        \timer_top_0/state_switch_0/N_293 ));
    NOR2B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m113  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[19] ), .B(
        \top_code_0_s_addchoice_5[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_114 ));
    AO1 \timer_top_0/state_switch_0/dataout_RNO[18]  (.A(
        \state_1ms_0_timecount[18] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .C(
        \timer_top_0/state_switch_0/N_270 ), .Y(
        \timer_top_0/state_switch_0/dataout_RNO[18]_net_1 ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[0]  (
        .D(\s_acq_change_0_s_acqnum[0] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load_0), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[0]_net_1 )
        );
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_97  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_153_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_70_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_18_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_97_Y ));
    DFN1 \PLUSE_0/qq_coder_0/i[0]  (.D(\PLUSE_0/qq_coder_0/i_RNO_7[0] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_9[0] ));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[9]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_177 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_178 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[9]_net_1 ));
    AX1 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m46  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i22_mux ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[12] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[13] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m46_4 ));
    DFN1 \PLUSE_0/qq_state_1/cs_i[0]  (.D(\PLUSE_0/qq_state_1/cs4 ), 
        .CLK(GLA_net_1), .Q(\PLUSE_0/qq_state_1/cs_i[0]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m142  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_135 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_142 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_143 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNI2E0P[13]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[13]_net_1 ), .B(
        \sd_acq_top_0/count_0[13] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_13[0] ));
    AND3 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_6_inst  
        (.A(\pd_pluse_top_0/count_6[3] ), .B(
        \pd_pluse_top_0/count_6[4] ), .C(\pd_pluse_top_0/count_1[5] ), 
        .Y(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_5_net ));
    NOR3A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[3]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/N_174 ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/N_175 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_0[3]_net_1 ));
    DFN1E1 \top_code_0/sigtimedata[0]  (.D(\GPMI_0_dataout[0] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[0] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_1[10]  (.A(
        \scanstate_0_timecount[10] ), .B(
        \timer_top_0/state_switch_0/N_295 ), .Y(
        \timer_top_0/state_switch_0/N_251 ));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_1_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ));
    OR3 \scalestate_0/timecount_ret_19_RNII8I  (.A(
        \scalestate_0/timecount_20_iv_3_reto[8] ), .B(
        \scalestate_0/timecount_20_iv_2_reto[8] ), .C(
        \scalestate_0/timecount_20_iv_6_reto[8] ), .Y(
        \scalestate_0/timecount_20_iv_9_reto[8] ));
    XOR2 \PLUSE_0/bri_timer_0/count_RNO[6]  (.A(
        \PLUSE_0/bri_timer_0/count_c5 ), .B(\PLUSE_0/count_2[6] ), .Y(
        \PLUSE_0/bri_timer_0/count_n6 ));
    DFN1E1 \state_1ms_0/PLUSETIME[10]  (.D(
        \top_code_0_state_1ms_data[10] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[10]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m268  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[14] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_269 ));
    AND3 \scalestate_0/necount_inc_0/AND2_5_inst  (.A(
        \scalestate_0/necount_inc_0/inc_2_net ), .B(
        \scalestate_0/necount[3]_net_1 ), .C(
        \scalestate_0/necount[4]_net_1 ), .Y(
        \scalestate_0/necount_inc_0/Rcout_5_net ));
    DFN1E1 \plusestate_0/timecount_1[7]  (.D(
        \plusestate_0/timecount_5[7] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[7] ));
    MX2 \state_1ms_0/timecount_RNO_0[18]  (.A(
        \state_1ms_0/timecount_8[18] ), .B(\state_1ms_0_timecount[18] )
        , .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_85 ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_22  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[2] ), .C(
        \timer_top_0/timer_0/DWACT_FINC_E[3] ), .Y(
        \timer_top_0/timer_0/N_15 ));
    DFN1 \timer_top_0/state_switch_0/dataout[20]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[20]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[20] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m25  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[8] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i14_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[8] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i16_mux ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_92  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_125_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_63_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_16_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_92_Y ));
    XOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf_RNIEF7R[0]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[0]_net_1 )
        , .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[0]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout8_0 ));
    DFN1E1 \top_code_0/plusedata[4]  (.D(\GPMI_0_dataout_0[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[4] ));
    DFN1E1 \state_1ms_0/M_DUMPTIME[14]  (.D(
        \top_code_0_state_1ms_data[14] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/M_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/M_DUMPTIME[14]_net_1 ));
    OA1 
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_0 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout14_NE_1 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/addrout[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ctrl_addr_0/addrout_RNIJIJB2[1]_net_1 )
        );
    AO1A \scalestate_0/timecount_ret_1_RNO_2  (.A(
        \scalestate_0/N_1089 ), .B(\scalestate_0/S_DUMPTIME[5]_net_1 ), 
        .C(\scalestate_0/timecount_20_iv_1[5] ), .Y(
        \scalestate_0/timecount_20_iv_6[5] ));
    OA1C \PLUSE_0/qq_state_0/cs_RNO_0[2]  (.A(Q3Q6_c), .B(
        \PLUSE_0/i_4[2] ), .C(\PLUSE_0/qq_state_0/cs[1]_net_1 ), .Y(
        \PLUSE_0/qq_state_0/N_89 ));
    DFN1E0 \DDS_0/dds_state_0/para[36]  (.D(
        \DDS_0/dds_state_0/para_9[36] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[36]_net_1 ));
    DFN1 \top_code_0/scale_rst_3  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_3));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[10]  (.D(
        \top_code_0_pd_pluse_data[10] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[10]_net_1 ));
    INV \GPMI_0/INV_0  (.A(gpio_c), .Y(\GPMI_0/INV_0_Y ));
    DFN1 \DUMP_ON_0/off_on_coder_0/i[1]  (.D(
        \DUMP_ON_0/off_on_coder_0/i_RNO_5[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_ON_0/i_5[1] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_122  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_73_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_21_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_15_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_122_Y ));
    AO1 \DUMP_0/dump_state_0/cs_RNI1C5R[7]  (.A(
        \DUMP_0/dump_state_0/un1_ns_0_a3_0 ), .B(
        \DUMP_0/dump_state_0/N_201 ), .C(
        \DUMP_0/dump_state_0/cs[7]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_168 ));
    DFN1 \timer_top_0/state_switch_0/dataout[4]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[4]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[4] ));
    AO1 \state_1ms_0/timecount_RNO_2[1]  (.A(
        \state_1ms_0/PLUSECYCLE[1]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[1] ), 
        .Y(\state_1ms_0/timecount_8_iv_1[1] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[9]  (.A(
        \plusestate_0_timecount[9] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_204 ));
    IOTRI_OR_EB \ddswclk_pad/U0/U1  (.D(
        \DDS_0/dds_state_0/w_clk_RNO_net_1 ), .E(VCC), .OCLK(GLA_net_1)
        , .DOUT(\ddswclk_pad/U0/NET1 ), .EOUT(\ddswclk_pad/U0/NET2 ));
    DFN1 \PLUSE_0/qq_coder_1/i[3]  (.D(\PLUSE_0/qq_coder_1/i_RNO_3[3] )
        , .CLK(GLA_net_1), .Q(\PLUSE_0/i_2[3] ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[0]  (.A(
        \top_code_0_dumpdata_0[0] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[0]_net_1 ));
    AO1A \DUMP_0/dump_state_0/timer_start_RNO_0  (.A(
        \DUMP_0/dump_state_0/N_168 ), .B(
        \DUMP_0/dump_state_0_timer_start ), .C(
        \DUMP_0/dump_state_0/ns[3] ), .Y(\DUMP_0/dump_state_0/N_88 ));
    DFN1E1 \top_code_0/pd_pluse_data[7]  (.D(\GPMI_0_dataout[7] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[7] ));
    AO1 \scalestate_0/timecount_ret_87_RNO  (.A(
        \scalestate_0/OPENTIME[10]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[10] ), .Y(
        \scalestate_0/timecount_20_iv_2[10] ));
    AO1 \scalestate_0/timecount_ret_8_RNO_2  (.A(
        \scalestate_0/CUTTIME180[3]_net_1 ), .B(\scalestate_0/N_263 ), 
        .C(\scalestate_0/OPENTIME_m[3] ), .Y(
        \scalestate_0/timecount_20_iv_2[3] ));
    DFN1E1 \top_code_0/change[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/change_1_sqmuxa ), .Q(
        \top_code_0_change[1] ));
    AO1 \state_1ms_0/timecount_RNO_2[14]  (.A(
        \state_1ms_0/M_DUMPTIME[14]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[14] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[14] ));
    AND2 \ClockManagement_0/clk_10k_0/un1_count_1_I_1  (.A(
        \ClockManagement_0/clk_10k_0/count[0]_net_1 ), .B(
        \ClockManagement_0/clk_5M_en ), .Y(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_TMP[0] ));
    NOR2A \scalestate_0/timecount_ret_77_RNO_4  (.A(
        \scalestate_0/CUTTIME90[6]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[6] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[18]  (.D(
        \top_code_0_sd_sacq_data[2] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_360 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[18]_net_1 ));
    NOR3C \DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa  (.A(
        \DUMP_OFF_1/off_on_state_0_state_over ), .B(
        nsctrl_choice_0_dumpoff_ctr), .C(nsctrl_choice_0_dumponoff_rst)
        , .Y(\DUMP_OFF_1/off_on_timer_0/count_0_sqmuxa_net_1 ));
    MX2 \scalestate_0/strippluse_RNO_0[0]  (.A(
        \scalestate_0/strippluse_6[0] ), .B(
        \scalestate_0_strippluse[0] ), .S(\scalestate_0/un1_CS6_26 ), 
        .Y(\scalestate_0/N_559 ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_4_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_4_net ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[3]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10_i ), .CLK(
        GLA_net_1), .E(top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall[3]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[13]_net_1 ));
    DFN1E1 \scanstate_0/timecount_1[0]  (.D(
        \scanstate_0/timecount_5[0] ), .CLK(GLA_net_1), .E(
        \scanstate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \scanstate_0_timecount[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/m46_3 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[13] ));
    NOR3C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO_0[11]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c10 ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[9]  (.A(
        \ClockManagement_0/long_timer_0/count_c8 ), .B(
        \ClockManagement_0/long_timer_0/count[9]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n9 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[11]  (.D(
        \top_code_0_sd_sacq_data[11] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[11]_net_1 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[16]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[16] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[16] ));
    NOR2B \nsctrl_choice_0/intertodsp_RNO  (.A(
        \nsctrl_choice_0/intertodsp_5 ), .B(net_27), .Y(
        \nsctrl_choice_0/intertodsp_RNO_net_1 ));
    DFN1E1 \top_code_0/sigtimedata[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[11] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m261  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[15] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_262 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i12_mux ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para1[2]  (.D(
        \top_code_0_bri_datain[2] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para1[2] ));
    XO1 \bridge_div_0/datahalf_RNIIC6F1[2]  (.A(
        \bridge_div_0/count[2]_net_1 ), .B(
        \bridge_div_0/datahalf[2]_net_1 ), .C(
        \bridge_div_0/clear1_n17_1[0] ), .Y(
        \bridge_div_0/clear1_n17_NE_1[0] ));
    OA1C \top_code_0/scanchoice_RNO  (.A(\top_code_0/N_208 ), .B(
        top_code_0_scanchoice), .C(\top_code_0/N_306 ), .Y(
        \top_code_0/N_98 ));
    DFN1E1 \top_code_0/bri_datain[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/bri_datain_1_sqmuxa ), .Q(
        \top_code_0_bri_datain[7] ));
    XOR3 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/un3_addresult_m69  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_2[1] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_4[1] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_2_i ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/N_70_i ));
    NOR2B \ClockManagement_0/long_timer_0/count_RNIJ5LR[5]  (.A(
        \ClockManagement_0/long_timer_0/count[5]_net_1 ), .B(
        \ClockManagement_0/long_timer_0/count[6]_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_m6_0_a2_2 ));
    XA1 \PLUSE_0/qq_timer_1/count_RNO[3]  (.A(
        \PLUSE_0/qq_timer_1/count_c2 ), .B(\PLUSE_0/count_7[3] ), .C(
        \PLUSE_0/qq_timer_1/count_0_sqmuxa_net_1 ), .Y(
        \PLUSE_0/qq_timer_1/count_n3 ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[15]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[15] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[15] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[5]  (.A(\s_acq_change_0/N_61 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[5]_net_1 ));
    MX2 \Signal_Noise_Acq_0/n_s_change_0/dataout[11]  (.A(
        \Signal_Noise_Acq_0/signal_data_t[11] ), .B(
        \Signal_Noise_Acq_0/MX2_RD_11_inst ), .S(top_code_0_n_s_ctrl_0)
        , .Y(\Signal_Noise_Acq_0_dataout[11] ));
    AOI1A \PLUSE_0/bri_coder_0/half_0_I_10  (.A(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[0] ), .B(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[1] ), .C(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[2] ), .Y(
        \PLUSE_0/bri_coder_0/ACT_LT3_E[3] ));
    NOR3B \top_code_0/scaledatain_1_sqmuxa_0_a2  (.A(
        \top_code_0/N_331 ), .B(\top_code_0/N_332 ), .C(
        \top_code_0/N_164 ), .Y(\top_code_0/scaledatain_1_sqmuxa ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_19[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[10]_net_1 ), 
        .B(\pd_pluse_top_0/count_0[10] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_10[0] ));
    AO1 \scalestate_0/timecount_ret_31_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL[4]_net_1 ), .B(
        \scalestate_0/N_261 ), .C(\scalestate_0/CUTTIME180_Tini_m[4] ), 
        .Y(\scalestate_0/timecount_20_iv_3[4] ));
    XOR2 \scalestate_0/M_pulse_RNO_12  (.A(
        \scalestate_0/M_NUM[0]_net_1 ), .B(
        \scalestate_0/necount[0]_net_1 ), .Y(\scalestate_0/M_pulse8_0 )
        );
    NOR2B \bridge_div_0/clk_4f_reg2_RNIREDC_0  (.A(
        \bridge_div_0/clk_4f_reg1_net_1 ), .B(
        \bridge_div_0/clk_4f_reg2_i_0 ), .Y(clk_4f_en_0));
    OR3 \scalestate_0/timecount_ret_37_RNI23EE  (.A(
        \scalestate_0/timecount_20_iv_7_reto[3] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[3] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[3] ), .Y(
        \scalestate_0/timecount_20_iv_10_reto[3] ));
    DFN1C0 \PLUSE_0/bri_coder_0/i[3]/U1  (.D(
        \PLUSE_0/bri_coder_0/i[3]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/i_3[3] ));
    DFN1E1 \top_code_0/n_divnum[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/n_divnum_1_sqmuxa ), .Q(
        \top_code_0_n_divnum_0[7] ));
    NOR2B \top_code_0/relay_on_RNO[7]  (.A(\top_code_0/N_816 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[7]_net_1 ));
    DFN1 \timer_top_0/state_switch_0/clk_en_st1ms  (.D(
        \timer_top_0/state_switch_0/clk_en_st1ms_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(timer_top_0_clk_en_st1ms));
    AO1A \DDS_0/dds_state_0/para_RNO_2[17]  (.A(
        \top_code_0_dds_configdata[0] ), .B(
        \DDS_0/dds_state_0/N_569_1 ), .C(\DDS_0/dds_state_0/N_498 ), 
        .Y(\DDS_0/dds_state_0/para_9_i_1[17] ));
    DFN1E1 \scalestate_0/timecount_ret_26  (.D(
        \scalestate_0/timecount_20_iv_8[11]_net_1 ), .CLK(GLA_net_1), 
        .E(\scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[11] ));
    OA1B \plusestate_0/CS_RNO[8]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[8]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[8] )
        , .Y(\plusestate_0/CS_RNO[8]_net_1 ));
    OR3 \top_code_0/nstatechoice_RNO_0  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_161 ), .Y(
        \top_code_0/N_210 ));
    DFN1E1 \top_code_0/dds_configdata[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[13] ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[5]  (.D(
        \DUMP_0/dump_coder_0/para2_4[5]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[5]_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_2[12]  (.A(
        \state_1ms_0/M_DUMPTIME[12]_net_1 ), .B(
        \state_1ms_0/CS[6]_net_1 ), .C(\state_1ms_0/PLUSECYCLE_m[12] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_0[12] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m130  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_129 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_130 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_131 ));
    DFN1E1 \bridge_div_0/dataall[1]  (.D(\bridge_div_0/dataall_1[1] ), 
        .CLK(GLA_net_1), .E(top_code_0_bridge_load), .Q(
        \bridge_div_0/dataall[1]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m181  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_178 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_181 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_182 ));
    OA1C \top_code_0/s_load_RNO  (.A(\top_code_0/N_196 ), .B(
        top_code_0_s_load), .C(\top_code_0/N_302 ), .Y(
        \top_code_0/N_94 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m61  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[5] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i8_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_62_i ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[13]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c12 ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[13]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n13 ));
    IOIN_IB \xa_pad[13]/U0/U1  (.YIN(\xa_pad[13]/U0/NET1 ), .Y(
        \xa_c[13] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m31  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i18_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[10] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i20_mux ));
    XA1C \sd_acq_top_0/sd_sacq_coder_0/i_RNO_5[10]  (.A(
        \sd_acq_top_0/count[18] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[18]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_3_14[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_3[10] ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[7]  (.D(
        \DUMP_0/dump_coder_0/para2_4[7]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[7]_net_1 ));
    NOR2B \top_code_0/relay_close_RNO[2]  (.A(\top_code_0/N_821 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[2]_net_1 ));
    NOR3C \scalestate_0/necount_LE_M_RNI0LLA  (.A(
        \scalestate_0/CS[15]_net_1 ), .B(
        \scalestate_0/necount_LE_M_net_1 ), .C(top_code_0_scale_rst_0), 
        .Y(\scalestate_0/N_261 ));
    MX2B \plusestate_0/timecount_1_RNO[0]  (.A(\plusestate_0/N_71 ), 
        .B(top_code_0_pluse_rst), .S(\plusestate_0/N_271 ), .Y(
        \plusestate_0/timecount_5[0] ));
    DFN1E1 \scalestate_0/timecount_ret_58  (.D(
        \scalestate_0/timecount_20_iv_6[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[0] ));
    AO1 \timer_top_0/timer_0/Timer_Cmp_0/AO1_2  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_5_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_4_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_0_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AO1_2_Y ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[9]  (.D(
        \top_code_0_pd_pluse_data[9] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[9]_net_1 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m109  (.A(
        \top_code_0_s_addchoice_1[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[4] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_110 ));
    IOPAD_TRI \relay_close_pad[2]/U0/U0  (.D(
        \relay_close_pad[2]/U0/NET1 ), .E(\relay_close_pad[2]/U0/NET2 )
        , .PAD(relay_close[2]));
    NOR2B \state_1ms_0/timecount_RNO_5[14]  (.A(
        \state_1ms_0/PLUSECYCLE[14]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[14] ));
    OA1B \noisestate_0/CS_RNO[7]  (.A(timer_top_0_clk_en_noise), .B(
        \noisestate_0/CS[7]_net_1 ), .C(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Y(
        \noisestate_0/CS_RNO[7]_net_1 ));
    DFN1 \state_1ms_0/pluse_start  (.D(\state_1ms_0/pluse_start_RNO_2 )
        , .CLK(GLA_net_1), .Q(state_1ms_0_pluse_start));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[3]  (.D(
        \top_code_0_pd_pluse_data[3] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[3]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[18]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[18]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_503 ));
    DFN1E0 \DUMP_0/dump_coder_0/para6[9]  (.D(
        \DUMP_0/dump_coder_0/para2_4[9]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para6[9]_net_1 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataseven[6]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataseven_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[6] ));
    DFN1E1 \scanstate_0/acqtime[1]  (.D(\top_code_0_scandata[1] ), 
        .CLK(GLA_net_1), .E(\scanstate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \scanstate_0/acqtime[1]_net_1 ));
    XOR2 \timer_top_0/timer_0/un2_timedata_I_28  (.A(
        \timer_top_0/timer_0/N_13 ), .B(
        \timer_top_0/timer_0/timedata[10]_net_1 ), .Y(
        \timer_top_0/timer_0/I_28_0 ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[6]  (.D(
        \top_code_0_scaledatain[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[6]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[6]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[7]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_277 ));
    DFN1E1 \plusestate_0/DUMPTIME[4]  (.D(\top_code_0_plusedata[4] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_1_sqmuxa_net_1 ), 
        .Q(\plusestate_0/DUMPTIME[4]_net_1 ));
    XA1A \timer_top_0/timer_0/Timer_Cmp_0/AND2_0  (.A(
        \timer_top_0/dataout[21] ), .B(
        \timer_top_0/timer_0/timedata[21]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_1_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND2_0_Y ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m19  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_12_0 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_19_0 ), .S(
        \top_code_0_s_addchoice_0[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_20 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNIIFJS[14]  (.A(
        \sd_acq_top_0/count_0[14] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[14]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_8[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_3[0] ));
    DFN1 \top_code_0/scale_rst_0_0  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_0));
    MX2 \top_code_0/noise_rst_0_0_RNIHP9S2  (.A(top_code_0_noise_rst_0)
        , .B(\xa_c[0] ), .S(\top_code_0/N_259 ), .Y(\top_code_0/N_805 )
        );
    DFN1 \DUMP_0/dump_state_0/cs[7]  (.D(
        \DUMP_0/dump_state_0/cs_nsss[7] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/dump_state_0/cs[7]_net_1 ));
    NOR2B \ClockManagement_0/clk_10k_0/clk_5M_reg1_RNO  (.A(net_27), 
        .B(\ClockManagement_0/pllclk_0_GLB ), .Y(
        \ClockManagement_0/clk_10k_0/clk_5M_reg1_RNO_net_1 ));
    DFN1 \timer_top_0/state_switch_0/dataout[9]  (.D(
        \timer_top_0/state_switch_0/dataout_RNO[9]_net_1 ), .CLK(
        GLA_net_1), .Q(\timer_top_0/dataout[9] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_1[1]  (.A(
        \top_code_0_s_acqnum_2[1] ), .B(\scalestate_0_s_acqnum[1] ), 
        .S(\top_code_0_change_0[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[1] ));
    NOR2B \scalestate_0/CS_RNIKC1B1[14]  (.A(\scalestate_0/N_1304 ), 
        .B(\scalestate_0/N_1266 ), .Y(\scalestate_0/N_1309 ));
    NOR2A \PLUSE_0/bri_state_0/cs_RNIB75I[11]  (.A(clk_4f_en), .B(
        \PLUSE_0/bri_state_0/cs[11]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/N_183 ));
    NOR2B \ClockManagement_0/long_timer_0/en  (.A(top_code_0_sigrst), 
        .B(net_27), .Y(\ClockManagement_0/long_timer_0/en_net_1 ));
    NOR2B \s_acq_change_0/s_acqnum_RNO[3]  (.A(\s_acq_change_0/N_73 ), 
        .B(net_27), .Y(\s_acq_change_0/s_acqnum_RNO[3]_net_1 ));
    AND2A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_44  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_52_i ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E[2] )
        );
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_2_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_17_Y ));
    DFN1E1 \scalestate_0/STRIPNUM90_NUM[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/STRIPNUM90_NUM_1_sqmuxa ), .Q(
        \scalestate_0/STRIPNUM90_NUM[5]_net_1 ));
    OR3 \state_1ms_0/timecount_RNO_1[0]  (.A(
        \state_1ms_0/timecount_8_0_iv_0[0] ), .B(
        \state_1ms_0/CUTTIME_m[0] ), .C(
        \state_1ms_0/timecount_8_0_iv_1[0] ), .Y(
        \state_1ms_0/timecount_8[0] ));
    XOR2 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_RNITKUE[5]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[5]_net_1 ), 
        .B(\pd_pluse_top_0/count_1[5] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_reg10_5[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[10]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[10]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_292 ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m70  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .B(
        \Signal_Noise_Acq_0/un1_n_s_change_0_1[0] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m70 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[3]_net_1 ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[1]  (.D(
        \top_code_0_pd_pluse_data[1] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[1]_net_1 ));
    NOR2A \scalestate_0/timecount_ret_65_RNO_4  (.A(
        \scalestate_0/CUTTIME90[13]_net_1 ), .B(\scalestate_0/N_1069 ), 
        .Y(\scalestate_0/CUTTIME90_m[13] ));
    NOR2A \top_code_0/pluse_str_RNO_3  (.A(\xa_c[7] ), .B(\xa_c[5] ), 
        .Y(\top_code_0/un1_xa_49_0_a2_1 ));
    NOR2B \s_acq_change_0/s_load_0_0_RNIEJ0I1  (.A(
        \s_acq_change_0/N_69 ), .B(net_27), .Y(
        \s_acq_change_0/s_load_0_0_RNIEJ0I1_net_1 ));
    OR3 \scalestate_0/timecount_ret_64_RNO  (.A(
        \scalestate_0/ACQTIME_m[13] ), .B(
        \scalestate_0/PLUSETIME90_m[13] ), .C(
        \scalestate_0/S_DUMPTIME_m[13] ), .Y(
        \scalestate_0/timecount_20_iv_6[13] ));
    NOR3B \scalestate_0/PLUSETIME90_0_sqmuxa_0_a2  (.A(
        \scalestate_0/N_61 ), .B(\scalestate_0/N_62 ), .C(
        \top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/PLUSETIME90_0_sqmuxa ));
    DFN1 \noisestate_0/CS[3]  (.D(\noisestate_0/CS_RNO[3]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[3]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[1]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_70_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[1] ));
    NOR2B \scalestate_0/strippluse_RNO[5]  (.A(\scalestate_0/N_564 ), 
        .B(top_code_0_scale_rst), .Y(
        \scalestate_0/strippluse_RNO[5]_net_1 ));
    OR3 \scalestate_0/timecount_ret_51_RNIA4I  (.A(
        \scalestate_0/timecount_20_0_iv_0_reto[18] ), .B(
        \scalestate_0/OPENTIME_TEL_m_reto[18] ), .C(
        \scalestate_0/timecount_20_0_iv_4_reto[18] ), .Y(
        \scalestate_0_timecount[18] ));
    MX2 \scalestate_0/s_acqnum_1_RNO_1[3]  (.A(\scalestate_0/N_451 ), 
        .B(\scalestate_0/ACQECHO_NUM[3]_net_1 ), .S(
        \scalestate_0/CS_0[11]_net_1 ), .Y(
        \scalestate_0/s_acqnum_7[3] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[5]  (.D(
        \top_code_0_sd_sacq_data[5] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_394 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6[5]_net_1 ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIA2SG[10]  (.A(
        \DUMP_0/dump_coder_0/para3[10]_net_1 ), .B(\DUMP_0/count[10] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_10[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m195  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_194 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_195 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_196 ));
    MX2 \top_code_0/pluse_rst_0_0_RNIS8853  (.A(top_code_0_pluse_rst_0)
        , .B(\xa_c[0] ), .S(\top_code_0/N_264 ), .Y(\top_code_0/N_804 )
        );
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_stripnum_I_29  
        (.A(\s_acq_change_0_s_stripnum[6] ), .B(
        \s_acq_change_0_s_stripnum[7] ), .C(
        \s_acq_change_0_s_stripnum[8] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_FINC_E[5] )
        );
    XOR2 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/XOR2_4_inst  (.A(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/Rcout_5_net ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[5] ));
    OR3 \scalestate_0/timecount_ret_58_RNO  (.A(
        \scalestate_0/ACQTIME_m[0] ), .B(
        \scalestate_0/PLUSETIME90_m[0] ), .C(
        \scalestate_0/S_DUMPTIME_m[0] ), .Y(
        \scalestate_0/timecount_20_iv_6[0] ));
    NOR2B \state_1ms_0/timecount_RNO_5[12]  (.A(
        \state_1ms_0/PLUSECYCLE[12]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .Y(\state_1ms_0/PLUSECYCLE_m[12] ));
    AOI1 \DUMP_OFF_1/off_on_state_0/cs_RNI1RQ6[1]  (.A(
        DUMP_OFF_1_dump_off), .B(\DUMP_OFF_1/i_4[1] ), .C(
        \DUMP_OFF_1/off_on_state_0/cs[1]_net_1 ), .Y(
        \DUMP_OFF_1/off_on_state_0/N_42_i ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_5[10]  (.A(
        \scalestate_0_timecount[10] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_253 ));
    OR2A \top_code_0/bri_datain_1_sqmuxa_0_o2  (.A(\xa_c[0] ), .B(
        \top_code_0/N_149 ), .Y(\top_code_0/N_160 ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/half_para[5]  (.D(
        \top_code_0_halfdata_0[5] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load), .Q(\PLUSE_0/half_para[5] ));
    IOTRI_OB_EB \sd_acq_en_pad/U0/U1  (.D(sd_acq_en_c), .E(VCC), .DOUT(
        \sd_acq_en_pad/U0/NET1 ), .EOUT(\sd_acq_en_pad/U0/NET2 ));
    OR3 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI07602[1]  (
        .A(\pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_0[0] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_4[0] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_7[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_11[0] ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_6  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/NOR3A_0_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_13_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_11_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_6_Y ));
    NOR3B \DUMP_0/dump_coder_0/i_RNO[7]  (.A(
        state1ms_choice_0_reset_out), .B(
        \DUMP_0/dump_coder_0/i_reg16_NE[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO[7]_net_1 ));
    NOR2B \scalestate_0/timecount_RNO_1[21]  (.A(
        \scalestate_0/OPENTIME_TEL[21]_net_1 ), .B(
        \scalestate_0/N_258 ), .Y(\scalestate_0/OPENTIME_TEL_m[21] ));
    MX2 \top_code_0/relay_close_RNO_0[0]  (.A(\relay_close_c[0] ), .B(
        \GPMI_0_dataout_0[0] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_819 ));
    NOR2B \scalestate_0/necount_RNO[4]  (.A(\scalestate_0/N_734 ), .B(
        top_code_0_scale_rst_4), .Y(
        \scalestate_0/necount_RNO[4]_net_1 ));
    MX2 \noisestate_0/timecount_1_RNO_0[4]  (.A(
        \noisestate_0/acqtime[4]_net_1 ), .B(
        \noisestate_0/dectime[4]_net_1 ), .S(\noisestate_0/N_191 ), .Y(
        \noisestate_0/N_61 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIEQ0P[19]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[19]_net_1 ), .B(
        \sd_acq_top_0/count[19] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_19[0] ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[11]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[11] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[11] ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_50_e  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_2_i_a2_0_net_1 )
        , .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_sd_sacq_data117_3_i_a2_1 ), 
        .C(\top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ));
    XOR2 \DSTimer_0/dump_sustain_timer_0/start_RNO_3  (.A(
        \DSTimer_0/dump_sustain_timer_0/data[1]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/count[1]_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/un1_data_1 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[16]  (.A(
        \scalestate_0_timecount[16] ), .B(
        \timer_top_0/state_switch_0/N_168 ), .Y(
        \timer_top_0/state_switch_0/N_266 ));
    DFN1E1 \state_1ms_0/PLUSETIME[9]  (.D(
        \top_code_0_state_1ms_data[9] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[9]_net_1 ));
    DFN1E1 \scalestate_0/PLUSETIME90[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME90_0_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME90[13]_net_1 ));
    AND3 \timer_top_0/timer_0/Timer_Cmp_0/AND3_2  (.A(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_3_Y ), .B(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_10_Y ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_18_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/AND3_2_Y ));
    AX1C \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m42  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[16] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_39_i ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[17] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/m42_4 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_7  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_7_Y ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[4]  (.A(\s_acq_change_0/N_60 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[4]_net_1 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_14_0  (.A(\xd_in[0] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout_0[0] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIC41I1[16]  (.A(
        \sd_acq_top_0/count[16] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[16]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_14[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_2[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[17]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_382 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[17]_net_1 ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_RNI5CD71[2]  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[0]_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[2] ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count_c2 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_3[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_3[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_64_i ));
    IOPAD_TRI \pd_pulse_en_pad/U0/U0  (.D(\pd_pulse_en_pad/U0/NET1 ), 
        .E(\pd_pulse_en_pad/U0/NET2 ), .PAD(pd_pulse_en));
    MX2 \plusestate_0/timecount_1_RNO_0[14]  (.A(
        \plusestate_0/PLUSETIME[14]_net_1 ), .B(
        \plusestate_0/DUMPTIME[14]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_85 ));
    DFN1E1 \state_1ms_0/PLUSETIME[15]  (.D(
        \top_code_0_state_1ms_data[15] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSETIME_1_sqmuxa ), .Q(
        \state_1ms_0/PLUSETIME[15]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_70  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_1_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_70_Y ));
    DFN1E1 \scalestate_0/ACQECHO_NUM[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ), .Q(
        \scalestate_0/ACQECHO_NUM[1]_net_1 ));
    DFN1E1 \top_code_0/scaledatain_0[1]  (.D(\GPMI_0_dataout_0[1] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain_0[1] ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_6  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_46_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[0] )
        );
    DFN1E1 \top_code_0/sd_sacq_data[1]  (.D(\GPMI_0_dataout[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[1] ));
    MX2 \plusestate_0/soft_d_RNO_0  (.A(\plusestate_0/N_302 ), .B(
        plusestate_0_soft_d), .S(\plusestate_0/N_299 ), .Y(
        \plusestate_0/N_121 ));
    DFN1 \bri_dump_sw_0/off_test  (.D(
        \bri_dump_sw_0/off_test_RNO_net_1 ), .CLK(GLA_net_1), .Q(
        bri_dump_sw_0_off_test));
    DFN1 \top_code_0/relay_close[4]  (.D(
        \top_code_0/relay_close_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_close_c[4] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m16  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[5] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i8_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[5] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i10_mux ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[13]  (.D(
        \top_code_0_sd_sacq_data[13] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[13]_net_1 ));
    DFN1 \noisestate_0/CS[2]  (.D(\noisestate_0/CS_RNO[2]_net_1 ), 
        .CLK(GLA_net_1), .Q(\noisestate_0/CS[2]_net_1 ));
    XNOR3 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/dataall_1_m9  (.A(
        \top_code_0_n_divnum_0[3] ), .B(\top_code_0_n_divnum_0[8] ), 
        .C(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/i4_mux ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/N_10_i ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m189  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_182 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_189 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[11] ));
    DFN1 \DUMP_OFF_0/off_on_timer_0/count[4]  (.D(
        \DUMP_OFF_0/off_on_timer_0/count_n4 ), .CLK(GLA_net_1), .Q(
        \DUMP_OFF_0/count_3[4] ));
    NOR2B \state_1ms_0/timecount_RNO_3[0]  (.A(
        \state_1ms_0/CUTTIME[0]_net_1 ), .B(\state_1ms_0/CS[8]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_m[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m150  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_147 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_150 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_151 ));
    DFN1E1 \top_code_0/pd_pluse_data[3]  (.D(\GPMI_0_dataout_0[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[19]  (
        .D(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/ADD_20x20_slow_I19_Y_1 )
        , .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[19] ));
    OA1B \state_1ms_0/CS_RNO[8]  (.A(\state_1ms_0/CS[8]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(\state_1ms_0/CS_srsts_i_0[8] ), 
        .Y(\state_1ms_0/CS_RNO_1[8] ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[0]  (.D(
        \DUMP_0/dump_coder_0/para5_4[0] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[0]_net_1 ));
    NOR2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[8] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_2_Y ));
    OR3A \scalestate_0/rt_sw_RNO_1  (.A(\scalestate_0/N_1195 ), .B(
        \scalestate_0/CS[13]_net_1 ), .C(\scalestate_0/N_1210 ), .Y(
        \scalestate_0/un1_CS_34 ));
    XNOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_5  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[10]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_44_i ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_1[1] )
        );
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[6]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n6 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ));
    AOI1A 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_34  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[3] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[6] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/ACT_LT4_E_0[10] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_CMPLE_PO0_DWACT_COMP0_E[2] )
        );
    OR2A \scalestate_0/necount_cmp_0/OR2A_2  (.A(
        \scalestate_0/M_NUM[8]_net_1 ), .B(
        \scalestate_0/necount[8]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_2_Y ));
    DFN1 \DUMP_0/off_on_state_0/cs[0]  (.D(
        \DUMP_0/off_on_state_0/N_36_i ), .CLK(GLA_net_1), .Q(
        DUMP_0_dump_off));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[7]  (.D(
        \top_code_0_sd_sacq_data[7] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[7]_net_1 ));
    DFN1 \sd_acq_top_0/sd_sacq_state_0/cs[5]  (.D(
        \sd_acq_top_0/sd_sacq_state_0/cs_RNO_3[5] ), .CLK(ddsclkout_c), 
        .Q(\sd_acq_top_0/sd_sacq_state_0/cs[5]_net_1 ));
    NOR2B \scalestate_0/timecount_ret_48_RNO_0  (.A(
        \scalestate_0/CUTTIME180[17]_net_1 ), .B(\scalestate_0/N_263 ), 
        .Y(\scalestate_0/CUTTIME180_m[17] ));
    OR3C \timer_top_0/timer_0/timedata_RNO[0]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/timedata[0]_net_1 ), .Y(
        \timer_top_0/timer_0/timedata_4[0] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORB_GATE_12_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/NOR2_0_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2_3_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEBP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_12_net ));
    NOR3A \DUMP_0/dump_state_0/cs_RNO[2]  (.A(
        \DUMP_0/dump_state_0/cs4 ), .B(\DUMP_0/dump_state_0/N_182 ), 
        .C(\DUMP_0/dump_state_0/N_183 ), .Y(
        \DUMP_0/dump_state_0/cs_RNO[2]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_Tini[16]  (.D(
        \top_code_0_scaledatain[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1745 ), .Q(
        \scalestate_0/CUTTIME180_Tini[16]_net_1 ));
    MX2B \noisestate_0/timecount_1_RNO[3]  (.A(\noisestate_0/N_60 ), 
        .B(\noisestate_0/N_193 ), .S(\noisestate_0/N_228 ), .Y(
        \noisestate_0/timecount_5[3] ));
    DFN1E1 \top_code_0/state_1ms_data[12]  (.D(\GPMI_0_dataout[12] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[12] ));
    RAM512X18 #( .MEMORYFILE("RAM_R6C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R6C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_6_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_6_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_0_net ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_115  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR10_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR11_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_115_Y ));
    NOR3B \DSTimer_0/dump_sustain_timer_0/start_RNO  (.A(
        \DSTimer_0/dump_sustain_timer_0/start11_0 ), .B(
        \DSTimer_0/dump_sustain_timer_0/start11_1 ), .C(
        \DSTimer_0/dump_sustain_timer_0/un1_data_0 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/start11 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[8]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_56_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[8] ));
    DFN1 \DUMP_0/off_on_state_0/cs[1]  (.D(
        \DUMP_0/off_on_state_0/cs_nsss[1] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/off_on_state_0/cs[1]_net_1 ));
    OA1 \top_code_0/un1_state_1ms_rst_n117_43_i_a3_0  (.A(
        \top_code_0/N_326 ), .B(\top_code_0/N_325 ), .C(
        \top_code_0/un1_state_1ms_rst_n117_43_i_a3_0_0_net_1 ), .Y(
        \top_code_0/N_328 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[1]  (.D(
        \top_code_0_scaledatain_0[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[1]_net_1 ));
    NOR2B \DUMP_ON_0/off_on_timer_0/count_RNO_0[4]  (.A(
        \DUMP_ON_0/count_5[3] ), .B(
        \DUMP_ON_0/off_on_timer_0/count_c2 ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_9_0 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[16]  (.A(
        \DDS_0/dds_state_0/N_535_0 ), .B(
        \DDS_0/dds_state_0/para_reg[16]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_296 ));
    DFN1 \top_code_0/relay_on[5]  (.D(
        \top_code_0/relay_on_RNO[5]_net_1 ), .CLK(GLA_net_1), .Q(
        \relay_on_c[5] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[10]  (.D(
        \top_code_0_sd_sacq_data[10] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[10]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[1]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIMEI90[18]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1767 ), .Q(\scalestate_0/CUTTIMEI90[18]_net_1 )
        );
    IOIN_IB \xa_pad[16]/U0/U1  (.YIN(\xa_pad[16]/U0/NET1 ), .Y(
        \xa_c[16] ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[9]  (.D(
        \ClockManagement_0/long_timer_0/count_n9 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[9]_net_1 ));
    NOR3B \bridge_div_0/count_RNIFNOM7[1]  (.A(pd_pulse_en_c), .B(
        \bridge_div_0/count[1]_net_1 ), .C(\bridge_div_0/clear1_n18 ), 
        .Y(\bridge_div_0/count_RNIFNOM7[1]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m49  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[11] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i20_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_50_i ));
    MX2 \PLUSE_0/bri_coder_0/i[4]/U0  (.A(\PLUSE_0/i_1[4] ), .B(
        bri_dump_sw_0_turn_delay), .S(clk_4f_en_0), .Y(
        \PLUSE_0/bri_coder_0/i[4]/Y ));
    DFN1E0 \DUMP_0/dump_coder_0/para1[10]  (.D(
        \DUMP_0/dump_coder_0/para4_4[10]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_6_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para1[10]_net_1 ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/un3_addresult_m41  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/N_41_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[18] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m41 ));
    OR2A \scalestate_0/necount_cmp_0/OR2A_5  (.A(
        \scalestate_0/necount[5]_net_1 ), .B(
        \scalestate_0/M_NUM[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_5_Y ));
    MX2B \scalestate_0/CS_RNO_0[1]  (.A(\scalestate_0/CS[1]_net_1 ), 
        .B(\scalestate_0/CS_i[0]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(\scalestate_0/N_1217 ));
    OA1C \top_code_0/pn_change_RNO  (.A(\top_code_0/N_219 ), .B(
        top_code_0_pn_change), .C(\top_code_0/N_300 ), .Y(
        \top_code_0/N_92 ));
    DFN1E1 \noisestate_0/timecount_1[7]  (.D(
        \noisestate_0/timecount_5[7] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[7] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[11]  (.A(
        \s_acq_change_0/s_acqnum_5[11] ), .B(
        \s_acq_change_0_s_acqnum[11] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_81 ));
    AND3 \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/AND2b_9_inst  (.A(
        \sd_acq_top_0/count_10[0] ), .B(\sd_acq_top_0/count_10[1] ), 
        .C(\sd_acq_top_0/count_10[2] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_2_net ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_1_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[3]_net_1 ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[5]  (.D(
        \top_code_0_scaledatain[5] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[5]_net_1 ));
    NOR2A \DUMP_0/dump_state_0/cs_RNO_1[4]  (.A(\DUMP_0/i_2[1] ), .B(
        \DUMP_0/dump_state_0/cs[4]_net_1 ), .Y(
        \DUMP_0/dump_state_0/N_186 ));
    DFN1E1 \state_1ms_0/CUTTIME[1]  (.D(\top_code_0_state_1ms_data[1] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[1]_net_1 ));
    NOR2A 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datafour_0  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        );
    DFN1 \s_acq_change_0/s_acqnum[12]  (.D(
        \s_acq_change_0/s_acqnum_RNO[12]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[12] ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m238  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[7] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_239 ));
    NOR3C \scalestate_0/timecount_ret_31_RNO_0  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[4]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[4] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_RD_1_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_130_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_139_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_0_Y ), .Y(
        \Signal_Noise_Acq_0/MX2_RD_1_inst ));
    DFN1 \DDS_0/dds_state_0/cs[4]  (.D(
        \DDS_0/dds_state_0/cs_RNO[4]_net_1 ), .CLK(GLA_net_1), .Q(
        \DDS_0/dds_state_0/cs[4]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_2/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_2/m46 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_6[13] ));
    NOR2B 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/en_net_1 ), .B(
        n_acq_change_0_n_rst_n), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        );
    DFN1 \pd_pluse_top_0/pd_pluse_state_0/stateover  (.D(
        \pd_pluse_top_0/pd_pluse_state_0/stateover_RNO_net_1 ), .CLK(
        ddsclkout_c), .Q(\pd_pluse_top_0/pd_pluse_state_0_stateover ));
    MX2A \noisestate_0/n_acq_RNO_0  (.A(\noisestate_0/N_191 ), .B(
        noisestate_0_n_acq), .S(\noisestate_0/N_229 ), .Y(
        \noisestate_0/N_129 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[32]  (.A(
        \DDS_0/dds_state_0/N_534 ), .B(
        \DDS_0/dds_state_0/para[33]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_314 ));
    DFN1E1 \top_code_0/sd_sacq_load  (.D(\top_code_0/N_102 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_sd_sacq_load));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[0]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m70_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[0] ));
    NOR3B \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk_RNO  (
        .A(top_code_0_n_rd_en), .B(n_acq_change_0_n_rst_n), .C(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/un1_clk_wire ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk_syn_0/n_rdclk_RNO_net_1 )
        );
    AO1B \scalestate_0/CS_RNIR1C72_0[18]  (.A(\scalestate_0/N_1310 ), 
        .B(timer_top_0_clk_en_scale_0), .C(top_code_0_scale_rst_0), .Y(
        \scalestate_0/un1_CS6_33_2 ));
    NOR2A \state_1ms_0/timecount_RNO_6[2]  (.A(
        \state_1ms_0/CS[8]_net_1 ), .B(\state_1ms_0/CUTTIME[2]_net_1 ), 
        .Y(\state_1ms_0/CUTTIME_i_m[2] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_23  (.A(
        \timer_top_0/dataout[16] ), .B(
        \timer_top_0/timer_0/timedata[16]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_23_Y ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNIVIQR8[10]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_14[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE_13[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_NE[0] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3_RNI9ET7[8]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data3[8]_net_1 ), .B(
        \sd_acq_top_0/count_1[8] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_5_8[0] ));
    OR2 \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_2[0]  (.A(
        \sd_acq_top_0/count[16] ), .B(\sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_19_2[0]_net_1 ));
    NOR2A \plusestate_0/timecount_1_RNO[13]  (.A(\plusestate_0/N_84 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[13] ));
    NOR2B \dds_change_0/dds_rst_RNO_2  (.A(net_45), .B(
        \top_code_0_change[0] ), .Y(\dds_change_0/ddsrstin2_m ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[10]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n10 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ));
    XO1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_RNI0K301[7]  (
        .A(\pd_pluse_top_0/count_1[7] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[7]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_5[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_NE_3[0] ));
    DFN1E1 \noisestate_0/acqtime[4]  (.D(\top_code_0_noisedata[4] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[4]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_57  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR6_11_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR7_11_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_57_Y ));
    XOR2 
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_1_5_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_7_net ), 
        .B(\pd_pluse_top_0/count_1[7] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[7] ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNISIO1[2]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c2 ));
    NOR2 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addrout[3] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addrout[2] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_dataone_2_net_1 )
        );
    OA1 \PLUSE_0/bri_coder_0/half_0_I_24  (.A(
        \PLUSE_0/bri_coder_0/N_11 ), .B(\PLUSE_0/bri_coder_0/N_10 ), 
        .C(\PLUSE_0/bri_coder_0/N_9 ), .Y(
        \PLUSE_0/bri_coder_0/DWACT_COMP0_E[2] ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_7_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_9_net ), 
        .B(\pd_pluse_top_0/count_0[9] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[9] ));
    DFN1 \top_code_0/scale_rst_5  (.D(
        \top_code_0/scale_rst_0_0_RNI25ID3_net_1 ), .CLK(GLA_net_1), 
        .Q(top_code_0_scale_rst_5));
    DFN1E1 \top_code_0/pd_pluse_data[2]  (.D(\GPMI_0_dataout_0[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[2] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]  (.D(
        \top_code_0_n_acqnum_2[8] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[8]_net_1 ));
    NOR3C \CAL_0/cal_div_0/count_RNO[3]  (.A(net_33_0), .B(
        \CAL_0/cal_div_0/cal_1_sqmuxa_1 ), .C(\CAL_0/cal_div_0/I_9 ), 
        .Y(\CAL_0/cal_div_0/count_5[3] ));
    OR2A \timer_top_0/timer_0/Timer_Cmp_0/OR2A_5  (.A(
        \timer_top_0/dataout[8] ), .B(
        \timer_top_0/timer_0/timedata[8]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_5_Y ));
    DFN1E1 \top_code_0/sd_sacq_data[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/sd_sacq_data_1_sqmuxa ), .Q(
        \top_code_0_sd_sacq_data[6] ));
    NOR3A \top_code_0/acqclken_RNO_1  (.A(\xa_c[2] ), .B(
        \top_code_0/N_151 ), .C(\top_code_0/N_165 ), .Y(
        \top_code_0/N_268 ));
    DFN1 \PLUSE_0/qq_state_0/cs_i[0]  (.D(\PLUSE_0/qq_state_0/cs4 ), 
        .CLK(GLA_net_1), .Q(\PLUSE_0/qq_state_0/cs_i[0]_net_1 ));
    NOR2B \DUMP_0/off_on_timer_0/count_RNIBU8J[2]  (.A(
        \DUMP_0/off_on_timer_0/count_c1 ), .B(\DUMP_0/count_2[2] ), .Y(
        \DUMP_0/off_on_timer_0/count_c2 ));
    DFN1E1 \top_code_0/sigrst  (.D(\top_code_0/N_104 ), .CLK(GLA_net_1)
        , .E(net_27), .Q(top_code_0_sigrst));
    DFN1 \plusestate_0/CS[8]  (.D(\plusestate_0/CS_RNO[8]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS[8]_net_1 ));
    DFN1E1 \top_code_0/dds_configdata[2]  (.D(\GPMI_0_dataout[2] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[2] ));
    DFN1C0 \GPMI_0/rst_n_module_0/rst_nr2  (.D(
        \GPMI_0/rst_n_module_0/rst_nr1_net_1 ), .CLK(GLA_net_1), .CLR(
        \GPMI_0/INV_0_Y ), .Q(\GPMI_0/rst_n_module_0/rst_nr2_net_1 ));
    AO1A \scalestate_0/timecount_ret_68_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[14]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[14] ), .Y(
        \scalestate_0/timecount_20_iv_0[14] ));
    DFN1E1 \top_code_0/scaledatain[13]  (.D(\GPMI_0_dataout[13] ), 
        .CLK(GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[13] ));
    DFN1E1 \scalestate_0/S_DUMPTIME[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[13]_net_1 ));
    DFN1C0 \GPMI_0/rst_n_module_0/rst_nr1  (.D(VCC), .CLK(GLA_net_1), 
        .CLR(\GPMI_0/INV_0_Y ), .Q(
        \GPMI_0/rst_n_module_0/rst_nr1_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_52  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_4_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_4_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_14_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_52_Y ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIP4PK[7]  (.A(
        \DUMP_0/dump_coder_0/para6[7]_net_1 ), .B(\DUMP_0/count_0[7] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_7[0] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_1[4]  (.A(
        \DDS_0/dds_state_0/N_535 ), .B(
        \DDS_0/dds_state_0/para_reg[4]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_317 ));
    DFN1E1 \top_code_0/dds_configdata[15]  (.D(\GPMI_0_dataout[15] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dds_configdata_1_sqmuxa ), .Q(
        \top_code_0_dds_configdata[15] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/un3_addresult_m59  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_5[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[6] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/i10_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_60_i ));
    OA1C \PLUSE_0/qq_state_0/cs_RNO_0[3]  (.A(
        \PLUSE_0/qq_state_0/cs[3]_net_1 ), .B(\PLUSE_0/i_4[3] ), .C(
        Q3Q6_c), .Y(\PLUSE_0/qq_state_0/N_86 ));
    NOR2A \GPMI_0/tri_state_0/dataout_1_3  (.A(\xd_in[11] ), .B(
        tri_ctrl_c), .Y(\GPMI_0_dataout[11] ));
    AO1 \DDS_0/dds_state_0/para_RNO[35]  (.A(
        \DDS_0/dds_state_0/para[35]_net_1 ), .B(
        \DDS_0/dds_state_0/N_538_1 ), .C(\DDS_0/dds_state_0/N_526 ), 
        .Y(\DDS_0/dds_state_0/para_9[35] ));
    NOR3 \PLUSE_0/bri_state_0/cs_RNO_9[3]  (.A(
        \PLUSE_0/bri_state_0/cs[8]_net_1 ), .B(
        \PLUSE_0/bri_state_0/cs[2]_net_1 ), .C(\PLUSE_0/i_3[2] ), .Y(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_7 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m231  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[8] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_232 ));
    DFN1E1 \scalestate_0/DUMPTIME[7]  (.D(\top_code_0_scaledatain[7] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/DUMPTIME[7]_net_1 ));
    XNOR2 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_22  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[6] ), 
        .B(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[6]_net_1 ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/DWACT_BL_EQUAL_0_E[2] )
        );
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/dataone[10]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[10] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_dataone ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0[10] ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[14]  
        (.D(\s_acq_change_0_s_acqnum[14] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[14]_net_1 )
        );
    DFN1 \timer_top_0/timer_0/timedata[6]  (.D(
        \timer_top_0/timer_0/timedata_4[6] ), .CLK(GLA_net_1), .Q(
        \timer_top_0/timer_0/timedata[6]_net_1 ));
    MX2B \state_1ms_0/pluse_start_RNO_0  (.A(state_1ms_0_pluse_start), 
        .B(\state_1ms_0/N_254 ), .S(\state_1ms_0/N_257 ), .Y(
        \state_1ms_0/N_155 ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m162  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[18] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_163 ));
    MX2B \topctrlchange_0/sw_acq1_RNO_0  (.A(sw_acq1_c), .B(
        \topctrlchange_0/sw_acq1_6_iv ), .S(
        \dds_change_0.un1_change_2 ), .Y(\topctrlchange_0/N_10 ));
    MX2 \state_1ms_0/timecount_RNO_0[4]  (.A(
        \state_1ms_0/timecount_8[4] ), .B(\state_1ms_0_timecount[4] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_71 ));
    DFN1E1 \noisestate_0/timecount_1[13]  (.D(
        \noisestate_0/timecount_5[13] ), .CLK(GLA_net_1), .E(
        \noisestate_0/un1_dumpoff_ctr_2_sqmuxa ), .Q(
        \noisestate_0_timecount[13] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n9 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[9]_net_1 )
        );
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr[7]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n7 ), .CLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .CLR(
        top_code_0_RAM_Rd_rst), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr[7] ));
    DFN1E1 \top_code_0/dump_cho[2]  (.D(\GPMI_0_dataout[2] ), .CLK(
        GLA_net_1), .E(\top_code_0/dump_cho_1_sqmuxa ), .Q(
        \top_code_0_dump_cho_0[2] ));
    DFN1E1 \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[3]  (.D(
        \top_code_0_n_divnum_0[3] ), .CLK(GLA_net_1), .E(
        top_code_0_n_load), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/datahalf[3]_net_1 ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_RNI8EKD[7]  (.A(
        \sd_acq_top_0/count_3[7] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2[7]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_5[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE_2[0] ));
    DFN1 \s_acq_change_0/s_acqnum[8]  (.D(
        \s_acq_change_0/s_acqnum_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_acqnum[8] ));
    NOR3C \scalestate_0/timecount_ret_64_RNO_1  (.A(
        top_code_0_scale_rst_3), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[13]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[13] ));
    XOR2 \DUMP_0/dump_coder_0/para6_RNIHSOK[3]  (.A(
        \DUMP_0/dump_coder_0/para6[3]_net_1 ), .B(\DUMP_0/count_1[3] ), 
        .Y(\DUMP_0/dump_coder_0/i_reg16_3[0] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult[4] ));
    XOR2 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m45  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_37_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[14] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m45_5 ));
    NOR2B \scalestate_0/rt_sw_RNO  (.A(\scalestate_0/N_544 ), .B(
        top_code_0_scale_rst_5), .Y(\scalestate_0/rt_sw_RNO_1_net_1 ));
    DFN1E0 \DDS_0/dds_state_0/para[8]  (.D(\DDS_0/dds_state_0/N_12 ), 
        .CLK(GLA_net_1), .E(\DDS_0/dds_state_0/para_1_sqmuxa_1 ), .Q(
        \DDS_0/dds_state_0/para[8]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[3]  (.D(\GPMI_0_dataout_0[3] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[3] ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[8]  (.A(
        \ClockManagement_0/long_timer_0/count_c7 ), .B(
        \ClockManagement_0/long_timer_0/count[8]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n8 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNIKV5R2[1]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_5[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_4[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_11[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_13[0] ));
    NOR2B \PLUSE_0/qq_timer_0/count_RNIDGIK[1]  (.A(
        \PLUSE_0/count_9[1] ), .B(\PLUSE_0/count_9[0] ), .Y(
        \PLUSE_0/qq_timer_0/count_c1 ));
    OR2 \PLUSE_0/bri_state_0/down_RNO  (.A(\PLUSE_0/bri_state_0/N_145 )
        , .B(\PLUSE_0/bri_state_0/cs[9]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/down32 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_4/addresult[18]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_4/m41_6 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_2[18] ));
    DFN1E1 \scalestate_0/ACQTIME[7]  (.D(\top_code_0_scaledatain[7] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[7]_net_1 ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m219  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_212 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_219 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[9] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[0]  (.A(
        \s_acq_change_0/s_acqnum_5[0] ), .B(
        \s_acq_change_0_s_acqnum[0] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_70 ));
    AO1A \DDS_0/dds_state_0/para_RNO_2[6]  (.A(
        \DDS_0/dds_state_0/para[6]_net_1 ), .B(
        \DDS_0/dds_state_0/N_569 ), .C(\DDS_0/dds_state_0/N_274 ), .Y(
        \DDS_0/dds_state_0/para_9_i_0_1[6] ));
    DFN1E1 \top_code_0/sigtimedata[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/sigtimedata_1_sqmuxa ), .Q(
        \top_code_0_sigtimedata[5] ));
    NOR2B \scan_scale_sw_0/s_start_RNO  (.A(\scan_scale_sw_0/N_26 ), 
        .B(net_27), .Y(\scan_scale_sw_0/s_start_RNO_net_1 ));
    DFN1E1 \top_code_0/dumpdata[6]  (.D(\GPMI_0_dataout[6] ), .CLK(
        GLA_net_1), .E(\top_code_0/dumpdata_1_sqmuxa ), .Q(
        \top_code_0_dumpdata_0[6] ));
    OR3 \scalestate_0/timecount_RNO[20]  (.A(
        \scalestate_0/timecount_20_0_iv_0[20] ), .B(
        \scalestate_0/OPENTIME_TEL_m[20] ), .C(
        \scalestate_0/timecount_20_0_iv_1[20] ), .Y(
        \scalestate_0/timecount_20[20] ));
    NOR2A \noisestate_0/timecount_1_RNO[12]  (.A(\noisestate_0/N_69 ), 
        .B(\noisestate_0/N_228 ), .Y(\noisestate_0/timecount_5[12] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m67  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[2] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[2] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/N_68_i ));
    DFN1 \scalestate_0/soft_d  (.D(\scalestate_0/soft_d_RNO_2 ), .CLK(
        GLA_net_1), .Q(scalestate_0_soft_d));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m38  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_38_i ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[15] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_39_i ));
    OR3 \DUMP_0/dump_coder_0/para3_RNIK9U52[2]  (.A(
        \DUMP_0/dump_coder_0/un1_count_2_3[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_2_4[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE_3[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_2_NE_7[0] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/un3_addresult_m57  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_1[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[7] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/i12_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_58_i ));
    NOR3C 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datasix[6]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_0_net_1 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/un2_datasix_1 )
        , .C(\Signal_Noise_Acq_0/un1_n_s_change_0_1[6] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_5[6] ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_13  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[0] ), .B(
        \timer_top_0/timer_0/timedata[3]_net_1 ), .C(
        \timer_top_0/timer_0/timedata[4]_net_1 ), .Y(
        \timer_top_0/timer_0/N_18 ));
    DFN1E1 \state_1ms_0/CUTTIME[0]  (.D(\top_code_0_state_1ms_data[0] )
        , .CLK(GLA_net_1), .E(\state_1ms_0/N_364 ), .Q(
        \state_1ms_0/CUTTIME[0]_net_1 ));
    MX2 \scanstate_0/timecount_1_RNO_0[0]  (.A(
        \scanstate_0/dectime[0]_net_1 ), .B(
        \scanstate_0/acqtime[0]_net_1 ), .S(\scanstate_0/CS[4]_net_1 ), 
        .Y(\scanstate_0/N_58 ));
    DFN1E1 \top_code_0/s_acqnum[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[9] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[12]  (.D(
        \top_code_0_sd_sacq_data[12] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_344 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4[12]_net_1 ));
    AO1A \state_1ms_0/timecount_RNO_2[5]  (.A(
        \state_1ms_0/PLUSECYCLE[5]_net_1 ), .B(
        \state_1ms_0/CS[4]_net_1 ), .C(\state_1ms_0/PLUSETIME_i_m[5] ), 
        .Y(\state_1ms_0/timecount_8_iv_1[5] ));
    NOR2B \top_code_0/relay_on_RNO[8]  (.A(\top_code_0/N_817 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[8]_net_1 ));
    NOR3B \ClockManagement_0/clk_10k_0/count_RNO[8]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/I_38_0 ), .C(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_10k_0/count_5[8] ));
    AO1C \plusestate_0/CS_RNO_0[3]  (.A(\plusestate_0/CS[8]_net_1 ), 
        .B(timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \plusestate_0/CS_srsts_i_0[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[5]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_62_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[5] ));
    DFN1E1 \plusestate_0/timecount_1[11]  (.D(
        \plusestate_0/timecount_5[11] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[11] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[11]  (.D(
        \top_code_0_pd_pluse_data[11] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data2[11]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[3]  (.D(
        \top_code_0_sd_sacq_data[3] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[3]_net_1 ));
    NOR2A \s_acq_change_0/s_acqnum_RNO_1[15]  (.A(
        \top_code_0_s_acqnum_2[15] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_acqnum_5[15] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m82  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_75 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_82 ), .S(
        \top_code_0_s_addchoice[3] ), .Y(
        \Signal_Noise_Acq_0/signal_data_t[6] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_27  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_131_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_72_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_8_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_27_Y ));
    DFN1E1 \scalestate_0/OPENTIME[13]  (.D(
        \top_code_0_scaledatain[13] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1665 ), .Q(\scalestate_0/OPENTIME[13]_net_1 ));
    DFN1C0 \PLUSE_0/bri_state_0/down/U1  (.D(
        \PLUSE_0/bri_state_0/down/Y ), .CLK(ddsclkout_c), .CLR(
        \PLUSE_0/bri_state_0/en_net_1 ), .Q(\PLUSE_0/down ));
    MX2 \scalestate_0/s_acqnum_1_RNO_0[4]  (.A(
        \scalestate_0/s_acqnum_7[4] ), .B(\scalestate_0_s_acqnum[4] ), 
        .S(\scalestate_0/un1_CS6_26 ), .Y(\scalestate_0/N_551 ));
    XOR2 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNO[7]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_c6 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n7 ));
    XOR2 \top_code_0/un1_state_1ms_rst_n117_28_i_o3  (.A(\xa_c[1] ), 
        .B(\xa_c[0] ), .Y(\top_code_0/N_169 ));
    NOR2B \top_code_0/relay_on_RNO[2]  (.A(\top_code_0/N_811 ), .B(
        net_27), .Y(\top_code_0/relay_on_RNO[2]_net_1 ));
    NOR3B 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_NE_7_RNISICAI6  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE ), 
        .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_i ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_65 ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ));
    NOR3A \PLUSE_0/qq_state_1/cs_RNO[3]  (.A(\PLUSE_0/qq_state_1/cs4 ), 
        .B(\PLUSE_0/qq_state_1/N_86 ), .C(\PLUSE_0/qq_state_1/N_87 ), 
        .Y(\PLUSE_0/qq_state_1/cs_RNO_2[3] ));
    DFN1E1 \scalestate_0/timecount_ret_77  (.D(
        \scalestate_0/timecount_20_iv_8[6] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[6] ));
    NOR3C \scalestate_0/timecount_ret_40_RNO_1  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[19]_net_1 ), .C(
        \scalestate_0/PLUSETIME90[2]_net_1 ), .Y(
        \scalestate_0/PLUSETIME90_m[2] ));
    NOR2B \topctrlchange_0/soft_dump_6_iv_RNO_0  (.A(
        plusestate_0_soft_d), .B(\top_code_0_change[1] ), .Y(
        \topctrlchange_0/s_dumpin3_m ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[11]  (.A(
        \plusestate_0_timecount[11] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_199 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m258  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[15] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_259 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[13]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/m46_5 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[13] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[1]  (.D(
        \top_code_0_sd_sacq_data[1] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_0_sqmuxa ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[1]_net_1 ));
    XOR2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_6_inst  
        (.A(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/Rcout_8_net ), 
        .B(\pd_pluse_top_0/count_0[8] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[8] ));
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[14]  (.D(
        \top_code_0_pd_pluse_data[14] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1_0_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data1[14]_net_1 ));
    NOR3 \DDS_0/dds_state_0/para_RNO[5]  (.A(\DDS_0/dds_state_0/N_323 )
        , .B(\DDS_0/dds_state_0/N_321 ), .C(
        \DDS_0/dds_state_0/para_9_i_1[5] ), .Y(
        \DDS_0/dds_state_0/N_81 ));
    IOBI_IB_OB_EB \xd_pad[10]/U0/U1  (.D(
        \Signal_Noise_Acq_0_dataout[10] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .YIN(\xd_pad[10]/U0/NET3 ), .DOUT(
        \xd_pad[10]/U0/NET1 ), .EOUT(\xd_pad[10]/U0/NET2 ), .Y(
        \xd_in[10] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_22  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_9_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_9_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_22_Y ));
    XO1 \DUMP_0/dump_coder_0/para5_RNIQCB71[2]  (.A(
        \DUMP_0/count_1[2] ), .B(\DUMP_0/dump_coder_0/para5[2]_net_1 ), 
        .C(\DUMP_0/dump_coder_0/un1_count_1_0[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE_3[0] ));
    OR3B \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ORA_GATE_5_inst  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_2_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/AND2A_0_Y ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/WEAP ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_5_net ));
    OA1B \plusestate_0/CS_RNO[9]  (.A(timer_top_0_clk_en_pluse), .B(
        \plusestate_0/CS[9]_net_1 ), .C(\plusestate_0/CS_srsts_i_0[9] )
        , .Y(\plusestate_0/CS_RNO[9]_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_timer_0/count_RNO[14]  (.A(
        pulse_start_c), .B(\pd_pluse_top_0/pd_pluse_state_0_stateover )
        , .C(\pd_pluse_top_0/pd_pluse_timer_0/count1[14] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[14] ));
    OR3 \DUMP_0/dump_coder_0/para2_RNI00SD2[0]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_10[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_3_0_0[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_3_NE_5[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_3_NE_8[0] ));
    XOR2 \DUMP_0/dump_coder_0/para5_RNIAJLJ[0]  (.A(
        \DUMP_0/dump_coder_0/para5[0]_net_1 ), .B(\DUMP_0/count_1[0] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_0[0] ));
    NOR3C \PLUSE_0/qq_coder_1/i_RNO[1]  (.A(
        \PLUSE_0/qq_coder_1/i_0_4[1] ), .B(
        \PLUSE_0/qq_coder_1/un1_qq_para2_i[0] ), .C(
        \PLUSE_0/qq_coder_1/i_reg10_NE[0]_net_1 ), .Y(
        \PLUSE_0/qq_coder_1/i_RNO_7[1] ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI3C3A[4]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[4]_net_1 ), .B(
        \sd_acq_top_0/count_10[4] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_4[0] ));
    AO1A \scalestate_0/timecount_20_iv_5_RNO[4]  (.A(
        \scalestate_0/N_1065 ), .B(\scalestate_0/ACQTIME[4]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[4] ), .Y(
        \scalestate_0/timecount_20_iv_0[4] ));
    DFN1E1 \scalestate_0/S_DUMPTIME[3]  (.D(
        \top_code_0_scaledatain_0[3] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[3]_net_1 ));
    AX1C \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/XOR2_3_inst  
        (.A(\pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_2_net )
        , .B(\pd_pluse_top_0/count_6[3] ), .C(
        \pd_pluse_top_0/count_6[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/count1[4] ));
    NOR2 \DUMP_0/dump_state_0/cs_srsts_0_0_a2_0[6]  (.A(\DUMP_0/i[7] ), 
        .B(\DUMP_0/i[5] ), .Y(\DUMP_0/dump_state_0/N_206 ));
    NOR2B \state_1ms_0/pluse_start_RNO  (.A(\state_1ms_0/N_155 ), .B(
        top_code_0_state_1ms_rst_n), .Y(
        \state_1ms_0/pluse_start_RNO_2 ));
    XOR2 \scalestate_0/M_pulse_RNO_13  (.A(
        \scalestate_0/M_NUM[2]_net_1 ), .B(
        \scalestate_0/necount[2]_net_1 ), .Y(\scalestate_0/M_pulse8_2 )
        );
    DFN1E1 \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[11]  (.D(
        \top_code_0_pd_pluse_data[11] ), .CLK(GLA_net_1), .E(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3_1_sqmuxa ), .Q(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[11]_net_1 ));
    DFN1E1 \top_code_0/s_acqnum[1]  (.D(\GPMI_0_dataout_0[1] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[1] ));
    XA1 \DUMP_ON_0/off_on_timer_0/count_RNO[4]  (.A(
        \DUMP_ON_0/off_on_timer_0/count_9_0 ), .B(
        \DUMP_ON_0/count_5[4] ), .C(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_n4 ));
    XA1 \DUMP_ON_0/off_on_timer_0/count_RNO[3]  (.A(
        \DUMP_ON_0/off_on_timer_0/count_c2 ), .B(
        \DUMP_ON_0/count_5[3] ), .C(
        \DUMP_ON_0/off_on_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DUMP_ON_0/off_on_timer_0/count_n3 ));
    AO1 \state_1ms_0/timecount_RNO_4[3]  (.A(
        \state_1ms_0/S_DUMPTIME[3]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CUTTIME_m[3] ), .Y(
        \state_1ms_0/timecount_8_iv_2[3] ));
    NOR3C \timer_top_0/timer_0/timedata_RNO[3]  (.A(net_27), .B(
        \timer_top_0/timer_0/time_up_0_sqmuxa_1 ), .C(
        \timer_top_0/timer_0/I_9_2 ), .Y(
        \timer_top_0/timer_0/timedata_4[3] ));
    DFN1E1 \scalestate_0/timecount_ret_23  (.D(
        \scalestate_0/timecount_20_iv_8[10] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[10] ));
    NOR2B \Signal_Noise_Acq_0/n_s_change_0/n_adc_1_4  (.A(\ADC_c[6] ), 
        .B(top_code_0_n_s_ctrl), .Y(\Signal_Noise_Acq_0/n_adc_1_4 ));
    DFN1 \scanstate_0/rt_sw  (.D(\scanstate_0/rt_sw_RNO_2 ), .CLK(
        GLA_net_1), .Q(scanstate_0_rt_sw));
    IOTRI_OB_EB \relay_on_pad[9]/U0/U1  (.D(\relay_on_c[9] ), .E(VCC), 
        .DOUT(\relay_on_pad[9]/U0/NET1 ), .EOUT(
        \relay_on_pad[9]/U0/NET2 ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_4  (.A(
        \timer_top_0/dataout[19] ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_4_Y ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[3]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_37 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[3] ));
    XOR2 \ClockManagement_0/clk_10k_0/un1_count_1_I_38  (.A(
        \ClockManagement_0/clk_10k_0/count[8]_net_1 ), .B(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_g_array_3[0] ), .Y(
        \ClockManagement_0/clk_10k_0/I_38_0 ));
    DFN1E1 \top_code_0/noisedata[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/noisedata_1_sqmuxa ), .Q(
        \top_code_0_noisedata[4] ));
    OR2 \scalestate_0/necount_LE_M_RNISD8P1  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_7_0 ), .B(
        \scalestate_0/N_263 ), .Y(
        \scalestate_0/un1_timecount_2_sqmuxa_7 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m296  (.A(
        \top_code_0_s_addchoice[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[12] ), .C(
        \top_code_0_s_addchoice_3[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_297 ));
    DFN1E1 \scalestate_0/S_DUMPTIME[15]  (.D(
        \top_code_0_scaledatain[15] ), .CLK(GLA_net_1), .E(
        \scalestate_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \scalestate_0/S_DUMPTIME[15]_net_1 ));
    AND2 \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/AND2_8_inst  
        (.A(\pd_pluse_top_0/count_1[6] ), .B(
        \pd_pluse_top_0/count_1[7] ), .Y(
        \pd_pluse_top_0/pd_pluse_timer_0/pd_pluse_inc_0/inc_8_net ));
    DFN1E1 \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[10]  
        (.D(\s_acq_change_0_s_acqnum[10] ), .CLK(GLA_net_1), .E(
        s_acq_change_0_s_load), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[10]_net_1 )
        );
    OR2A \scalestate_0/CS_RNI62781_0[17]  (.A(\scalestate_0/N_1194 ), 
        .B(\scalestate_0/N_1265 ), .Y(\scalestate_0/N_1209_0 ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[6]  (.A(
        \s_acq_change_0/s_acqnum_5[6] ), .B(
        \s_acq_change_0_s_acqnum[6] ), .S(\top_code_0_change_0[1] ), 
        .Y(\s_acq_change_0/N_76 ));
    NOR2B \scanstate_0/CS_i_0_RNI7I3Q[0]  (.A(\scanstate_0/CS_li[0] ), 
        .B(\scanstate_0/N_255 ), .Y(\scanstate_0/N_253 ));
    DFN1E1 \top_code_0/s_acqnum[5]  (.D(\GPMI_0_dataout[5] ), .CLK(
        GLA_net_1), .E(\top_code_0/s_acqnum_1_sqmuxa ), .Q(
        \top_code_0_s_acqnum_2[5] ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m22  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[7] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i12_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[7] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i14_mux ));
    NOR3B \scalestate_0/ACQECHO_NUM_1_sqmuxa_0_a2  (.A(
        \scalestate_0/N_60 ), .B(\scalestate_0/N_67 ), .C(
        \top_code_0_scalechoice_0_0[0] ), .Y(
        \scalestate_0/ACQECHO_NUM_1_sqmuxa ));
    MX2 \top_code_0/relay_close_RNO_0[5]  (.A(\relay_close_c[5] ), .B(
        \GPMI_0_dataout[5] ), .S(\top_code_0/relay_close_1_sqmuxa ), 
        .Y(\top_code_0/N_824 ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m251  (.A(
        \top_code_0_s_addchoice_4[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[15] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_252 ));
    DFN1 \DUMP_0/dump_timer_0/count[11]  (.D(
        \DUMP_0/dump_timer_0/count_n11 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count[11] ));
    DFN1 \top_code_0/inv_turn  (.D(\top_code_0/inv_turn_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(top_code_0_inv_turn));
    DFN1E1 \top_code_0/nstatechoice  (.D(\top_code_0/N_78 ), .CLK(
        GLA_net_1), .E(net_27), .Q(top_code_0_nstatechoice));
    MX2 \scalestate_0/pluse_start_RNO_0  (.A(\scalestate_0/N_1197 ), 
        .B(scalestate_0_pluse_start), .S(\scalestate_0/N_1171 ), .Y(
        \scalestate_0/N_725 ));
    NOR3C \DUMP_0/dump_timer_0/count_RNO_0[11]  (.A(\DUMP_0/count[9] ), 
        .B(\DUMP_0/dump_timer_0/count_c8 ), .C(
        \DUMP_0/dump_timer_0/count_23_0 ), .Y(
        \DUMP_0/dump_timer_0/N_52 ));
    OR3 \DUMP_0/dump_coder_0/para5_RNIOKBN7[0]  (.A(
        \DUMP_0/dump_coder_0/un1_count_NE_7[0] ), .B(
        \DUMP_0/dump_coder_0/un1_count_NE_6[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_NE_8[0] ), .Y(
        \DUMP_0/dump_coder_0/un1_count_NE[0] ));
    OA1A \PLUSE_0/bri_coder_0/half_0_I_19  (.A(\PLUSE_0/half_para[3] ), 
        .B(\PLUSE_0/count_8[3] ), .C(\PLUSE_0/bri_coder_0/N_3 ), .Y(
        \PLUSE_0/bri_coder_0/N_7 ));
    DFN1 \DUMP_0/dump_coder_0/i[0]  (.D(
        \DUMP_0/dump_coder_0/i_RNO_0[0] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_2[0] ));
    XNOR2 \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_20  (.A(
        \timer_top_0/dataout[19] ), .B(
        \timer_top_0/timer_0/timedata[19]_net_1 ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/XNOR2_20_Y ));
    RAM512X18 #( .MEMORYFILE("RAM_R9C0.mem") )  
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/RAM_R9C0  (.RADDR8(
        AFLSDF_GND), .RADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr[7] ), 
        .RADDR6(\Signal_Noise_Acq_0/noise_acq_0/addr[6] ), .RADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr[5] ), .RADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr[4] ), .RADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr[3] ), .RADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr[2] ), .RADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr[1] ), .RADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr[0] ), .WADDR8(AFLSDF_GND), 
        .WADDR7(\Signal_Noise_Acq_0/noise_acq_0/addr_0[7] ), .WADDR6(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .WADDR5(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .WADDR4(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[4] ), .WADDR3(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ), .WADDR2(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[2] ), .WADDR1(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[1] ), .WADDR0(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[0] ), .WD17(GND), .WD16(
        GND), .WD15(GND), .WD14(GND), .WD13(GND), .WD12(GND), .WD11(
        \Signal_Noise_Acq_0/n_adc_1 ), .WD10(
        \Signal_Noise_Acq_0/n_adc_1_0 ), .WD9(
        \Signal_Noise_Acq_0/n_adc_1_1 ), .WD8(
        \Signal_Noise_Acq_0/n_adc_1_2 ), .WD7(
        \Signal_Noise_Acq_0/n_adc_1_3 ), .WD6(
        \Signal_Noise_Acq_0/n_adc_1_4 ), .WD5(
        \Signal_Noise_Acq_0/n_adc_1_5 ), .WD4(
        \Signal_Noise_Acq_0/n_adc_1_6 ), .WD3(
        \Signal_Noise_Acq_0/n_adc_1_7 ), .WD2(
        \Signal_Noise_Acq_0/n_adc_1_8 ), .WD1(
        \Signal_Noise_Acq_0/n_adc_1_9 ), .WD0(
        \Signal_Noise_Acq_0/n_adc_1_10 ), .RW0(GND), .RW1(VCC), .WW0(
        GND), .WW1(VCC), .PIPE(GND), .REN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKB_EN_9_net ), .WEN(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BLKA_EN_9_net ), .RCLK(
        \Signal_Noise_Acq_0/noise_acq_0/n_rdclk ), .WCLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .RESET(
        n_acq_change_0_n_rst_n_0), .RD17(), .RD16(), .RD15(), .RD14(), 
        .RD13(), .RD12(), .RD11(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_11_net ), 
        .RD10(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_10_net ), 
        .RD9(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_9_net ), 
        .RD8(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_8_net ), 
        .RD7(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_7_net ), 
        .RD6(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_6_net ), 
        .RD5(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_5_net ), 
        .RD4(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_4_net ), 
        .RD3(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_3_net ), 
        .RD2(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_2_net ), 
        .RD1(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_1_net ), 
        .RD0(\Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_0_net ));
    DFN1C0 \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7]/U1  
        (.D(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7]/Y )
        , .CLK(\Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[7] ));
    XO1 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNILNRE1[7]  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[7]_net_1 )
        , .B(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/I_20 ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_6 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_6 ));
    NOR2B \sd_acq_top_0/sd_sacq_coder_0/i_RNO[3]  (.A(
        scalestate_0_long_opentime), .B(net_27), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_4[3] ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_44  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_16_Y ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_86_Y ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_10_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_44_Y ));
    NOR3B \DUMP_0/dump_coder_0/i_RNO[5]  (.A(
        \DUMP_0/dump_coder_0/N_19 ), .B(
        \DUMP_0/dump_coder_0/un1_count_1_NE[0] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/i_RNO[5]_net_1 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m63  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[4] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[4] ), 
        .C(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i6_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_64_i ));
    IOTRI_OB_EB \k1_pad/U0/U1  (.D(k1_c), .E(VCC), .DOUT(
        \k1_pad/U0/NET1 ), .EOUT(\k1_pad/U0/NET2 ));
    DFN1E1 \scalestate_0/timecount_ret_40  (.D(
        \scalestate_0/timecount_20_iv_6[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_1 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[2] ));
    DFN1E1 \scalestate_0/CUTTIME180[2]  (.D(
        \top_code_0_scaledatain_0[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1645 ), .Q(\scalestate_0/CUTTIME180[2]_net_1 ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/un3_addresult_m19  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult_0[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i10_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_6[6] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/i12_mux ));
    AX1C \ClockManagement_0/clk_div500_0/un1_count_1_I_37  (.A(
        \ClockManagement_0/clk_div500_0/DWACT_ADD_CI_0_g_array_1[0] ), 
        .B(\ClockManagement_0/clk_div500_0/count[2]_net_1 ), .C(
        \ClockManagement_0/clk_div500_0/count[3]_net_1 ), .Y(
        \ClockManagement_0/clk_div500_0/I_37 ));
    DFN1E1 \scalestate_0/timecount_ret_72  (.D(
        \scalestate_0/timecount_20_iv_6[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_6_reto[7] ));
    AOI1 \DUMP_0/off_on_state_1/cs_RNIIO2G[1]  (.A(DUMP_0_dump_on), .B(
        \DUMP_0/i_0[1] ), .C(\DUMP_0/off_on_state_1/cs[1]_net_1 ), .Y(
        \DUMP_0/off_on_state_1/N_42_i ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_0/addresult[4]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_0/N_64_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_5[4] ));
    DFN1C0 \pd_pluse_top_0/pd_pluse_timer_0/count[2]  (.D(
        \pd_pluse_top_0/pd_pluse_timer_0/count_3[2] ), .CLK(
        ddsclkout_c), .CLR(net_27), .Q(\pd_pluse_top_0/count_6[2] ));
    DFN1E1 \scalestate_0/CUTTIMEI90[11]  (.D(
        \top_code_0_scaledatain[11] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1751 ), .Q(\scalestate_0/CUTTIMEI90[11]_net_1 )
        );
    NOR2B \top_code_0/relay_close_RNO[4]  (.A(\top_code_0/N_823 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[4]_net_1 ));
    AX1C \sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/YXOR2_14_inst  (
        .A(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/incb_17_net ), 
        .B(\sd_acq_top_0/sd_sacq_timer_0/sd_sacq_inc_0/inc_28_net ), 
        .C(\sd_acq_top_0/count[18] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count1[18] ));
    OA1 \PLUSE_0/bri_state_0/cs_RNIVBIV[4]  (.A(\PLUSE_0/i_3[2] ), .B(
        \PLUSE_0/i_8[1] ), .C(\PLUSE_0/bri_state_0/cs[4]_net_1 ), .Y(
        \PLUSE_0/bri_state_0/N_181 ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data4_RNIGI6M3[3]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_1[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_0[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_NE_16[0] ));
    NOR2B \s_acq_change_0/s_stripnum_RNO_1[10]  (.A(
        \scalestate_0_strippluse[10] ), .B(\top_code_0_change[0] ), .Y(
        \s_acq_change_0/s_stripnum_5[10] ));
    MX2B \noisestate_0/timecount_1_RNO[9]  (.A(\noisestate_0/N_66 ), 
        .B(\noisestate_0/N_193 ), .S(\noisestate_0/N_228 ), .Y(
        \noisestate_0/timecount_5[9] ));
    OR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_RNI0GRB3[7]  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_8 )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_10 ), 
        .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_6 ), 
        .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk6_NE_10 )
        );
    DFN1 \scanstate_0/dds_conf  (.D(\scanstate_0/dds_conf_RNO_1 ), 
        .CLK(GLA_net_1), .Q(scanstate_0_dds_conf));
    NOR2B \DUMP_0/off_on_timer_1/count_RNO_0[4]  (.A(
        \DUMP_0/count_0[3] ), .B(\DUMP_0/off_on_timer_1/count_c2 ), .Y(
        \DUMP_0/off_on_timer_1/count_9_0 ));
    NOR2B \scalestate_0/timecount_ret_60_RNO_1  (.A(
        \scalestate_0/OPENTIME[12]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[12] ));
    OAI1 \scalestate_0/CS_RNO_0[8]  (.A(timer_top_0_clk_en_scale), .B(
        \scalestate_0/CS[8]_net_1 ), .C(top_code_0_scale_rst_3), .Y(
        \scalestate_0/CS_srsts_i_0[8] ));
    DFN1E1 \top_code_0/pd_pluse_data[0]  (.D(\GPMI_0_dataout_0[0] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[0] ));
    OR3 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data6_RNISU3S2[20]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_1[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_0[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_10[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_2_NE_16[0] ));
    OR2 \scalestate_0/CS_RNIVSUB[5]  (.A(\scalestate_0/CS[5]_net_1 ), 
        .B(\scalestate_0/CS[11]_net_1 ), .Y(\scalestate_0/N_1210 ));
    NOR2B 
        \Signal_Noise_Acq_0/signal_acq_0/ten_choice_one_0/datathree[9]  
        (.A(\Signal_Noise_Acq_0/un1_n_s_change_0_1[9] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/un2_datathree ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_2[9] ));
    NOR3C \scalestate_0/timecount_20_iv_5_RNO_1[11]  (.A(
        top_code_0_scale_rst_2), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[11]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[11] ));
    NOR2A \DDS_0/dds_state_0/cs_RNO[7]  (.A(\DDS_0/dds_state_0/N_223 ), 
        .B(\DDS_0/dds_state_0/N_226 ), .Y(\DDS_0/dds_state_0/N_80 ));
    DFN1E1 \CAL_0/cal_load_0/cal_para_out[2]  (.D(
        \top_code_0_cal_data[2] ), .CLK(GLA_net_1), .E(
        top_code_0_cal_load), .Q(\CAL_0/cal_para_out[2] ));
    DFN1E1 \PLUSE_0/bri_qq_load_0/qq_para3[2]  (.D(
        \top_code_0_bri_datain[12] ), .CLK(GLA_net_1), .E(
        top_code_0_bridge_load_0), .Q(\PLUSE_0/qq_para3[2] ));
    NOR3C 
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_RNIQF44[6]  
        (.A(\Signal_Noise_Acq_0/noise_acq_0/addr_0[5] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c4 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[6] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_c6 ));
    NOR2A \noisestate_0/CS_RNIRL68_0[1]  (.A(top_code_0_noise_rst), .B(
        \noisestate_0/CS[1]_net_1 ), .Y(
        \noisestate_0/timecount_cnst[2] ));
    NOR3C \scalestate_0/timecount_ret_38_RNO_3  (.A(
        top_code_0_scale_rst_1), .B(\scalestate_0/CS[20]_net_1 ), .C(
        \scalestate_0/PLUSETIME180[3]_net_1 ), .Y(
        \scalestate_0/PLUSETIME180_m[3] ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[2]  (.A(
        \top_code_0_dumpdata_0[2] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[2]_net_1 ));
    DFN1E1 \scalestate_0/M_NUM[0]  (.D(\top_code_0_scaledatain_0[0] ), 
        .CLK(GLA_net_1), .E(\scalestate_0/M_NUM_1_sqmuxa ), .Q(
        \scalestate_0/M_NUM[0]_net_1 ));
    DFN1E1 \top_code_0/n_rd_en  (.D(\top_code_0/N_74 ), .CLK(GLA_net_1)
        , .E(net_27), .Q(top_code_0_n_rd_en));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m198  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[10] ), .C(
        \top_code_0_s_addchoice_1[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_199 ));
    DFN1E1 \scalestate_0/ACQTIME[13]  (.D(\top_code_0_scaledatain[13] )
        , .CLK(GLA_net_1), .E(\scalestate_0/ACQTIME_1_sqmuxa ), .Q(
        \scalestate_0/ACQTIME[13]_net_1 ));
    NOR3C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_3[4]  (.A(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_2[4] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_1[4] ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_10[4] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_13[4] ));
    AO1 \state_1ms_0/timecount_RNO_4[10]  (.A(
        \state_1ms_0/S_DUMPTIME[10]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/PLUSETIME_m[10] ), 
        .Y(\state_1ms_0/timecount_8_0_iv_1[10] ));
    DFN1 \DUMP_0/dump_timer_0/count[5]  (.D(
        \DUMP_0/dump_timer_0/count_n5 ), .CLK(GLA_net_1), .Q(
        \DUMP_0/count_0[5] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]  (.D(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n6 ), 
        .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[6]_net_1 )
        );
    NOR2B \scalestate_0/timecount_ret_38_RNO_4  (.A(
        \scalestate_0/CUTTIMEI90[3]_net_1 ), .B(\scalestate_0/N_252 ), 
        .Y(\scalestate_0/CUTTIMEI90_m[3] ));
    NOR2B \DDS_0/dds_timer_0/count_RNI3HB8[0]  (.A(\DDS_0/count[0] ), 
        .B(\DDS_0/count[1] ), .Y(\DDS_0/dds_timer_0/count_c1 ));
    AO1A \scalestate_0/timecount_ret_71_RNO_0  (.A(
        \scalestate_0/N_1093 ), .B(\scalestate_0/DUMPTIME[15]_net_1 ), 
        .C(\scalestate_0/PLUSETIME180_m[15] ), .Y(
        \scalestate_0/timecount_20_iv_0[15] ));
    DFN1 \DUMP_0/dump_coder_0/i[2]  (.D(
        \DUMP_0/dump_coder_0/i_RNO_0[2] ), .CLK(GLA_net_1), .Q(
        \DUMP_0/i_0[2] ));
    NOR3B \timer_top_0/state_switch_0/state_start5_0_0_a2_1  (.A(
        \timer_top_0/state_switch_0/N_284 ), .B(
        \timer_top_0/state_switch_0/state_start5_0_0_a2_1_0_net_1 ), 
        .C(top_code_0_scale_start), .Y(
        \timer_top_0/state_switch_0/N_295 ));
    NOR2A \pd_pluse_top_0/pd_pluse_state_0/cs_RNO_1[3]  (.A(
        \pd_pluse_top_0/i_1[3] ), .B(
        \pd_pluse_top_0/pd_pluse_state_0/cs[2]_net_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/N_175 ));
    AO1C \state_1ms_0/CS_RNO_0[3]  (.A(\state_1ms_0/CS[2]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(\state_1ms_0/CS_srsts_i_0[3] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/addresult[14]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_1/m45_2 ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_4[14] ));
    OA1B \scanstate_0/CS_RNO[2]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[2]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[2] ), 
        .Y(\scanstate_0/CS_RNO_2[2] ));
    AO1A \scalestate_0/timecount_ret_4_RNIK9SS  (.A(
        \scalestate_0/un1_timecount_2_sqmuxa_reto ), .B(
        \scalestate_0/timecount_cnst_m_0_reto[2] ), .C(
        \scalestate_0/timecount_20_iv_10_reto[2] ), .Y(
        \scalestate_0_timecount[2] ));
    NOR2B \DDS_0/dds_timer_0/count_RNO_1[7]  (.A(\DDS_0/count[6] ), .B(
        \DDS_0/dds_timer_0/count_0_sqmuxa_net_1 ), .Y(
        \DDS_0/dds_timer_0/count_15_0 ));
    OA1C \top_code_0/dds_choice_RNO  (.A(\top_code_0/N_205 ), .B(
        top_code_0_dds_choice), .C(\top_code_0/N_274 ), .Y(
        \top_code_0/N_66 ));
    DFN1E1 \noisestate_0/acqtime[2]  (.D(\top_code_0_noisedata[2] ), 
        .CLK(GLA_net_1), .E(\noisestate_0/acqtime_1_sqmuxa_net_1 ), .Q(
        \noisestate_0/acqtime[2]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180[16]  (.D(
        \top_code_0_scaledatain_0[0] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1661 ), .Q(\scalestate_0/CUTTIME180[16]_net_1 )
        );
    NOR2A \DUMP_0/dump_coder_0/para2_4[2]  (.A(
        \top_code_0_dumpdata_0[2] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[2]_net_1 ));
    DFN1 \state_1ms_0/timecount[19]  (.D(
        \state_1ms_0/timecount_RNO[19]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[19] ));
    NOR2B \scalestate_0/timecount_ret_29_RNO_1  (.A(
        \scalestate_0/OPENTIME_TEL[1]_net_1 ), .B(\scalestate_0/N_258 )
        , .Y(\scalestate_0/OPENTIME_TEL_m[1] ));
    NOR3B \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_RNO[1]  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_0_sqmuxa_1_0_net_1 )
        , .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_5_1 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/clkout9 ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count_6[1] ));
    NOR2B \scalestate_0/dump_start_RNO  (.A(\scalestate_0/N_723 ), .B(
        top_code_0_scale_rst_5), .Y(
        \scalestate_0/dump_start_RNO_0_net_1 ));
    AO1 \scalestate_0/timecount_ret_71_RNO_2  (.A(
        \scalestate_0/CUTTIMEI90[15]_net_1 ), .B(\scalestate_0/N_252 ), 
        .C(\scalestate_0/CUTTIME90_m[15] ), .Y(
        \scalestate_0/timecount_20_iv_4[15] ));
    DFN1E1 \scalestate_0/OPENTIME_TEL[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1773 ), .Q(
        \scalestate_0/OPENTIME_TEL[7]_net_1 ));
    DFN1 \scalestate_0/sw_acq1  (.D(\scalestate_0/sw_acq1_RNO_0_net_1 )
        , .CLK(GLA_net_1), .Q(scalestate_0_sw_acq1));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m214  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_213 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_214 ), .S(
        \top_code_0_s_addchoice_1[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_215 ));
    NOR3C \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[7]  (.A(
        \pd_pluse_top_0/pd_pluse_state_0/en2 ), .B(
        \pd_pluse_top_0/i_0[4] ), .C(
        \pd_pluse_top_0/pd_pluse_state_0/cs_1 ), .Y(
        \pd_pluse_top_0/pd_pluse_state_0/cs_RNO[7]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_6/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_6/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_0[2] ));
    NOR3B \top_code_0/state_1ms_start_ret_2_RNO  (.A(
        \top_code_0/N_336 ), .B(\top_code_0/un1_xa_4_0_a2_1 ), .C(
        \top_code_0/N_163 ), .Y(\top_code_0/un1_xa_4 ));
    OA1B \scanstate_0/CS_RNO[3]  (.A(timer_top_0_clk_en_scan), .B(
        \scanstate_0/CS[3]_net_1 ), .C(\scanstate_0/CS_srsts_i_0[3] ), 
        .Y(\scanstate_0/CS_RNO_2[3] ));
    NOR2A \DUMP_0/dump_coder_0/para2_4[6]  (.A(
        \top_code_0_dumpdata_0[6] ), .B(\top_code_0_dump_cho_0[1] ), 
        .Y(\DUMP_0/dump_coder_0/para2_4[6]_net_1 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_167  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR2_10_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR3_10_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_6_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_167_Y ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/un3_count_I_12  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[3]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/DWACT_FINC_E[0] )
        , .C(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/count[4]_net_1 ), 
        .Y(\Signal_Noise_Acq_0/noise_acq_0/noiseclk_0/I_12_1 ));
    DFN1E1 \scalestate_0/timecount_ret_35  (.D(
        \scalestate_0/timecount_20_iv_8[9] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_0 ), .Q(
        \scalestate_0/timecount_20_iv_8_reto[9] ));
    MX2 \plusestate_0/timecount_1_RNO_0[6]  (.A(
        \plusestate_0/PLUSETIME[6]_net_1 ), .B(
        \plusestate_0/DUMPTIME[6]_net_1 ), .S(
        \plusestate_0/CS[5]_net_1 ), .Y(\plusestate_0/N_77 ));
    DFN1 \state_1ms_0/CS[6]  (.D(\state_1ms_0/CS_RNO_3[6] ), .CLK(
        GLA_net_1), .Q(\state_1ms_0/CS[6]_net_1 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_0[12]  (.A(
        \DDS_0/dds_state_0/N_534_0 ), .B(
        \DDS_0/dds_state_0/para[13]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_333 ));
    OR3 \scalestate_0/timecount_ret_14_RNI9SH  (.A(
        \scalestate_0/timecount_20_iv_7_reto[9] ), .B(
        \scalestate_0/timecount_20_iv_6_reto[9] ), .C(
        \scalestate_0/timecount_20_iv_8_reto[9] ), .Y(
        \scalestate_0/timecount_20_iv_10_reto[9] ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[28]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[28]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_478 ));
    OR2A 
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/un1_count_0_I_34  
        (.A(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/data[1]_net_1 ), 
        .B(\Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/count[1] ), 
        .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noiseclkctrl_0/ACT_LT4_E[1] ));
    OA1 \scalestate_0/CS_RNI0F0B[14]  (.A(\scalestate_0/CS[19]_net_1 ), 
        .B(\scalestate_0/CS[14]_net_1 ), .C(top_code_0_scale_rst_1), 
        .Y(\scalestate_0/un1_timecount_2_sqmuxa_6_1 ));
    DFN1C0 \sd_acq_top_0/sd_sacq_timer_0/count[19]  (.D(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[19] ), .CLK(ddsclkout_c), 
        .CLR(net_27), .Q(\sd_acq_top_0/count[19] ));
    OR3 \scalestate_0/timecount_ret_88_RNO  (.A(
        \scalestate_0/PLUSETIME90_m[10] ), .B(
        \scalestate_0/DUMPTIME_m[10] ), .C(
        \scalestate_0/S_DUMPTIME_m[10] ), .Y(
        \scalestate_0/timecount_20_iv_6[10] ));
    NOR3C \sd_acq_top_0/sd_sacq_timer_0/count_RNO[20]  (.A(
        scalestate_0_s_acq), .B(
        \sd_acq_top_0/sd_sacq_state_0_stateover ), .C(
        \sd_acq_top_0/sd_sacq_timer_0/count1[20] ), .Y(
        \sd_acq_top_0/sd_sacq_timer_0/count_3[20] ));
    NOR3B \scalestate_0/ACQTIME_1_sqmuxa_0_a2  (.A(\scalestate_0/N_60 )
        , .B(\scalestate_0/N_65 ), .C(\top_code_0_scalechoice_0_0[0] ), 
        .Y(\scalestate_0/ACQTIME_1_sqmuxa ));
    MX2 \bri_dump_sw_0/tetw_pluse_RNO_0  (.A(plusestate_0_tetw_pluse), 
        .B(scalestate_0_tetw_pluse), .S(top_code_0_pluse_scale), .Y(
        \bri_dump_sw_0/tetw_pluse_5 ));
    NOR2A \state_1ms_0/un1_PLUSECYCLE13_i_a2_0  (.A(
        top_code_0_state_1ms_load), .B(\top_code_0_state_1ms_lc[3] ), 
        .Y(\state_1ms_0/N_16 ));
    NOR2A \plusestate_0/timecount_1_RNO[15]  (.A(\plusestate_0/N_86 ), 
        .B(\plusestate_0/N_271 ), .Y(\plusestate_0/timecount_5[15] ));
    DFN1E1 \scalestate_0/timecount_ret_5  (.D(
        \scalestate_0/timecount_20_iv_7[2] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[2] ));
    AOI1B 
        \DSTimer_0/dump_sustain_timer_0/cmp_constant_4b_0/NAND2_AEB_RNIVFTG  
        (.A(\DSTimer_0/dump_sustain_timer_0/count[3]_net_1 ), .B(
        \DSTimer_0/dump_sustain_timer_0/cmp_constant_4b_0/Temp_0_net ), 
        .C(\DSTimer_0/dump_sustain_timer_0/enable_net_1 ), .Y(
        \DSTimer_0/dump_sustain_timer_0/un1_clr_cnt_p ));
    AO1A \top_code_0/noise_start_ret_3_RNO  (.A(\top_code_0/N_171 ), 
        .B(\top_code_0/un1_state_1ms_rst_n117_44_i_a2_0 ), .C(
        \top_code_0/N_162 ), .Y(\top_code_0/N_114 ));
    DFN1E1 \state_1ms_0/PLUSECYCLE[8]  (.D(
        \top_code_0_state_1ms_data[8] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/PLUSECYCLE_0_sqmuxa ), .Q(
        \state_1ms_0/PLUSECYCLE[8]_net_1 ));
    XOR2 \bridge_div_0/datahalf_RNI63JN[0]  (.A(
        \bridge_div_0/datahalf[0]_net_1 ), .B(
        \bridge_div_0/count[0]_net_1 ), .Y(
        \bridge_div_0/clear1_n17_0[0] ));
    NOR3A \top_code_0/pd_pluse_choice_1_sqmuxa_0_a2  (.A(
        \top_code_0/sigtimedata_1_sqmuxa_1 ), .B(\top_code_0/N_150 ), 
        .C(\top_code_0/N_167 ), .Y(
        \top_code_0/pd_pluse_choice_1_sqmuxa ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m51  
        (.A(\s_acq_change_0_s_stripnum[6] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[6]_net_1 )
        , .C(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i10_mux )
        , .Y(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_52_i ));
    XA1C \pd_pluse_top_0/pd_pluse_coder_0/i_RNO_7[4]  (.A(
        \pd_pluse_top_0/count_1[6] ), .B(
        \pd_pluse_top_0/pd_pluse_coder_0/pd_pluse_data3[6]_net_1 ), .C(
        \pd_pluse_top_0/pd_pluse_coder_0/un1_count_1_4[0] ), .Y(
        \pd_pluse_top_0/pd_pluse_coder_0/i_0_6[4] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[15]  (.A(
        \state_1ms_0_timecount[15] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_187 ));
    DFN1E1 \top_code_0/dump_sustain_data[3]  (.D(\GPMI_0_dataout[3] ), 
        .CLK(GLA_net_1), .E(\top_code_0/dump_sustain_data_1_sqmuxa ), 
        .Q(\top_code_0_dump_sustain_data[3] ));
    NAND3A \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_10  (.A(
        \timer_top_0/dataout[1] ), .B(
        \timer_top_0/timer_0/timedata[1]_net_1 ), .C(
        \timer_top_0/timer_0/Timer_Cmp_0/OR2A_2_Y ), .Y(
        \timer_top_0/timer_0/Timer_Cmp_0/NAND3A_10_Y ));
    OR2A \scalestate_0/necount_cmp_0/OR2A_0  (.A(
        \scalestate_0/M_NUM[5]_net_1 ), .B(
        \scalestate_0/necount[5]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/OR2A_0_Y ));
    NOR2A \PLUSE_0/qq_state_0/cs_RNII4451[4]  (.A(
        \PLUSE_0/qq_state_0/N_79 ), .B(
        \PLUSE_0/qq_state_0/cs[4]_net_1 ), .Y(
        \PLUSE_0/qq_state_0/N_84 ));
    NOR2A \DDS_0/dds_state_0/para_RNO_3[20]  (.A(
        \DDS_0/dds_state_0/N_538_1 ), .B(
        \DDS_0/dds_state_0/para[20]_net_1 ), .Y(
        \DDS_0/dds_state_0/N_466 ));
    DFN1E1 \scalestate_0/timecount_ret_60  (.D(
        \scalestate_0/timecount_20_iv_7[12] ), .CLK(GLA_net_1), .E(
        \scalestate_0/un1_CS6_33_2 ), .Q(
        \scalestate_0/timecount_20_iv_7_reto[12] ));
    DFN1E1 \top_code_0/plusedata[9]  (.D(\GPMI_0_dataout[9] ), .CLK(
        GLA_net_1), .E(\top_code_0/plusedata_1_sqmuxa ), .Q(
        \top_code_0_plusedata[9] ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_3/addresult[2]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_3/N_68_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_3[2] ));
    XOR2 \DUMP_0/dump_coder_0/para2_RNIFICG[4]  (.A(
        \DUMP_0/dump_coder_0/para2[4]_net_1 ), .B(\DUMP_0/count_1[4] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_3_4[0] ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[15]  (.D(
        \top_code_0_sd_sacq_data[15] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_410 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data7[15]_net_1 ));
    NOR3B \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa_0_a2  (
        .A(\sd_acq_top_0/sd_sacq_coder_0/N_24 ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/N_23 ), .C(
        \top_code_0_sd_sacq_choice[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data2_1_sqmuxa ));
    NOR2B \scalestate_0/timecount_ret_1_RNO_4  (.A(
        \scalestate_0/OPENTIME[5]_net_1 ), .B(\scalestate_0/N_259 ), 
        .Y(\scalestate_0/OPENTIME_m[5] ));
    DFN1 \ClockManagement_0/long_timer_0/clk_5K_reg1  (.D(
        \ClockManagement_0/long_timer_0/clk_5K_reg1_RNO_net_1 ), .CLK(
        GLA_net_1), .Q(
        \ClockManagement_0/long_timer_0/clk_5K_reg1_net_1 ));
    OR3A \ClockManagement_0/clk_10k_0/count_RNO[0]  (.A(net_27), .B(
        \ClockManagement_0/clk_10k_0/count_0_sqmuxa ), .C(
        \ClockManagement_0/clk_10k_0/DWACT_ADD_CI_0_partial_sum[0] ), 
        .Y(\ClockManagement_0/clk_10k_0/count_5[0] ));
    DFN1E1 \top_code_0/s_addchoice_4[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/s_addchoice_1_sqmuxa ), .Q(
        \top_code_0_s_addchoice_4[4] ));
    DFN1E1 \top_code_0/pd_pluse_data[11]  (.D(\GPMI_0_dataout[11] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[11] ));
    OR3 \timer_top_0/state_switch_0/dataout_RNO_2[13]  (.A(
        \timer_top_0/state_switch_0/N_192 ), .B(
        \timer_top_0/state_switch_0/N_194 ), .C(
        \timer_top_0/state_switch_0/N_193 ), .Y(
        \timer_top_0/state_switch_0/dataout_0_0_0_1[13] ));
    XO1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1_RNI24EB[4]  (.A(
        \sd_acq_top_0/count_10[4] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data1[4]_net_1 ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_6[0] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE_4[0] ));
    MX2 \top_code_0/scale_start_ret_RNIU5AM  (.A(
        \top_code_0/top_code_0_scale_start_reto ), .B(
        \top_code_0/xa_c_reto[0] ), .S(\top_code_0/N_110_reto ), .Y(
        \top_code_0/N_797_reto ));
    AO18 \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/un3_addresult_m34  
        (.A(\Signal_Noise_Acq_0/signal_acq_0/addresult[11] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i20_mux ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_7[11] ), 
        .Y(\Signal_Noise_Acq_0/signal_acq_0/add_reg_7/i22_mux ));
    AO1 \scalestate_0/timecount_ret_2_RNO_1  (.A(
        \scalestate_0/OPENTIME[6]_net_1 ), .B(\scalestate_0/N_259 ), 
        .C(\scalestate_0/CUTTIME180_m[6] ), .Y(
        \scalestate_0/timecount_20_iv_2[6] ));
    DFN1 \plusestate_0/CS_i[0]  (.D(\plusestate_0/CS_i_RNO[0]_net_1 ), 
        .CLK(GLA_net_1), .Q(\plusestate_0/CS_i[0]_net_1 ));
    DFN0C0 \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr[3]  (.D(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_0/addr_n3 ), .CLK(
        \Signal_Noise_Acq_0/s_clk_div4_0_clkout ), .CLR(
        n_acq_change_0_n_rst_n), .Q(
        \Signal_Noise_Acq_0/noise_acq_0/addr_0[3] ));
    MX2 \noisestate_0/timecount_1_RNO[5]  (.A(\noisestate_0/N_62 ), .B(
        top_code_0_noise_rst_0), .S(\noisestate_0/N_228 ), .Y(
        \noisestate_0/timecount_5[5] ));
    XA1 \ClockManagement_0/long_timer_0/count_RNO[6]  (.A(
        \ClockManagement_0/long_timer_0/count_c5 ), .B(
        \ClockManagement_0/long_timer_0/count[6]_net_1 ), .C(
        \ClockManagement_0/long_timer_0/en_net_1 ), .Y(
        \ClockManagement_0/long_timer_0/count_n6 ));
    NOR3A \scalestate_0/necount_cmp_0/NOR3A_1  (.A(
        \scalestate_0/necount_cmp_0/OR2A_2_Y ), .B(
        \scalestate_0/necount_cmp_0/AO1C_1_Y ), .C(
        \scalestate_0/M_NUM[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/NOR3A_1_Y ));
    AND3 \timer_top_0/timer_0/un2_timedata_I_45  (.A(
        \timer_top_0/timer_0/DWACT_FINC_E[6] ), .B(
        \timer_top_0/timer_0/DWACT_FINC_E[10] ), .C(
        \timer_top_0/timer_0/timedata[15]_net_1 ), .Y(
        \timer_top_0/timer_0/N_7 ));
    DFN1E1 \top_code_0/scaledatain[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/scaledatain_1_sqmuxa ), .Q(
        \top_code_0_scaledatain[7] ));
    NOR3B \ClockManagement_0/clk_div500_0/count_RNO[2]  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0/I_35 ), .C(
        \ClockManagement_0/clk_div500_0/count_0_sqmuxa ), .Y(
        \ClockManagement_0/clk_div500_0/count_5[2] ));
    MX2 \s_acq_change_0/s_acqnum_RNO_0[12]  (.A(
        \s_acq_change_0/s_acqnum_5[12] ), .B(
        \s_acq_change_0_s_acqnum[12] ), .S(\top_code_0_change[1] ), .Y(
        \s_acq_change_0/N_82 ));
    NOR2B \scalestate_0/s_acqnum_1_RNO[2]  (.A(\scalestate_0/N_549 ), 
        .B(top_code_0_scale_rst_5), .Y(
        \scalestate_0/s_acqnum_1_RNO[2]_net_1 ));
    AO1 \state_1ms_0/timecount_RNO_4[1]  (.A(
        \state_1ms_0/S_DUMPTIME[1]_net_1 ), .B(
        \state_1ms_0/CS[7]_net_1 ), .C(\state_1ms_0/CUTTIME_m[1] ), .Y(
        \state_1ms_0/timecount_8_iv_2[1] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m171  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_170 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_171 ), .S(
        \top_code_0_s_addchoice_2[0] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_172 ));
    XOR2 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5_RNI5E3A[5]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[5]_net_1 ), .B(
        \sd_acq_top_0/count_3[5] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_1_5[0] ));
    DFN1 \s_acq_change_0/s_stripnum[7]  (.D(
        \s_acq_change_0/s_stripnum_RNO[7]_net_1 ), .CLK(GLA_net_1), .Q(
        \s_acq_change_0_s_stripnum[7] ));
    DFN1E0C0 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count_n12 )
        , .CLK(\Signal_Noise_Acq_0/signal_acq_0/clkout ), .CLR(
        s_acq_change_0_s_rst), .E(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/enclk8 ), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/count[12]_net_1 )
        );
    IOTRI_OB_EB \Acq_clk_pad/U0/U1  (.D(Acq_clk_c), .E(VCC), .DOUT(
        \Acq_clk_pad/U0/NET1 ), .EOUT(\Acq_clk_pad/U0/NET2 ));
    NOR3C \DUMP_0/dump_coder_0/i_RNO_0[3]  (.A(
        \DUMP_0/dump_coder_0/un1_count_3_i[0] ), .B(
        \DUMP_0/dump_coder_0/i_0_0_a2_10[3] ), .C(
        \DUMP_0/dump_coder_0/un1_count_2_NE[0] ), .Y(
        \DUMP_0/dump_coder_0/i_0_0_a2_12[3] ));
    OR3 \scalestate_0/timecount_ret_14_RNO  (.A(
        \scalestate_0/CUTTIME180_TEL_m[9] ), .B(
        \scalestate_0/CUTTIME180_Tini_m[9] ), .C(
        \scalestate_0/timecount_20_iv_2[9] ), .Y(
        \scalestate_0/timecount_20_iv_7[9] ));
    NOR3C \PLUSE_0/qq_coder_1/i_RNO_0[1]  (.A(bri_dump_sw_0_reset_out), 
        .B(\PLUSE_0/qq_coder_1/i_0_1[1] ), .C(
        \PLUSE_0/qq_coder_1/i_0_2[1] ), .Y(
        \PLUSE_0/qq_coder_1/i_0_4[1] ));
    NOR2A \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m132  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[3] ), .B(
        \top_code_0_s_addchoice[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_133 ));
    AO1C \scalestate_0/necount_cmp_0/AO1C_1  (.A(
        \scalestate_0/necount[7]_net_1 ), .B(
        \scalestate_0/M_NUM[7]_net_1 ), .C(
        \scalestate_0/necount[6]_net_1 ), .Y(
        \scalestate_0/necount_cmp_0/AO1C_1_Y ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[0]  (.D(
        \ClockManagement_0/long_timer_0/N_95 ), .CLK(GLA_net_1), .E(
        \ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[0]_net_1 ));
    DFN1E1 \top_code_0/halfdata[7]  (.D(\GPMI_0_dataout[7] ), .CLK(
        GLA_net_1), .E(\top_code_0/halfdata_1_sqmuxa ), .Q(
        \top_code_0_halfdata_0[7] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_0[5]  (.A(
        \noisestate_0_timecount[5] ), .B(
        \timer_top_0/state_switch_0/N_296 ), .Y(
        \timer_top_0/state_switch_0/N_215 ));
    NOR3 \syn_md_module_1/syn_md_0/syn_md_out_RNO_1  (.A(
        \syn_md_module_1/syn_md_0/N_18 ), .B(
        \syn_md_module_1/syn_md_0/count[3]_net_1 ), .C(
        \syn_md_module_1/syn_md_edge_detect_0_syn_md_out_en ), .Y(
        \syn_md_module_1/syn_md_0/N_31 ));
    DFN1 \scalestate_0/s_acq  (.D(\scalestate_0/s_acq_RNO_net_1 ), 
        .CLK(GLA_net_1), .Q(scalestate_0_s_acq));
    BUFF \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/ADDRB_FF2_0_net ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_7_Y ));
    NOR2B \ClockManagement_0/long_timer_0/clk_5K_reg1_RNO  (.A(net_27), 
        .B(\ClockManagement_0/clk_div500_0_clk_5K ), .Y(
        \ClockManagement_0/long_timer_0/clk_5K_reg1_RNO_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para2[0]  (.D(
        \DUMP_0/dump_coder_0/para2_4[0]_net_1 ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_5_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para2[0]_net_1 ));
    IOPAD_TRI \sigtimeup_pad/U0/U0  (.D(\sigtimeup_pad/U0/NET1 ), .E(
        \sigtimeup_pad/U0/NET2 ), .PAD(sigtimeup));
    AND3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_count_1_0_I_8  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E_0[3] )
        , .B(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[4] )
        , .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_E[5] )
        , .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] )
        );
    NOR2A \scalestate_0/timecount_ret_58_RNO_0  (.A(
        \scalestate_0/ACQTIME[0]_net_1 ), .B(\scalestate_0/N_1065 ), 
        .Y(\scalestate_0/ACQTIME_m[0] ));
    NOR2A \scalestate_0/timecount_ret_33_RNI43C  (.A(
        \scalestate_0/timecount_m1_e_2_2_reto ), .B(
        \scalestate_0/un1_timecount_2_sqmuxa_9_reto ), .Y(
        \scalestate_0/timecount_cnst_m_reto[1] ));
    DFN1E1 \state_1ms_0/S_DUMPTIME[4]  (.D(
        \top_code_0_state_1ms_data[4] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/S_DUMPTIME_1_sqmuxa ), .Q(
        \state_1ms_0/S_DUMPTIME[4]_net_1 ));
    AO1 \PLUSE_0/bri_state_0/cs_RNO[3]  (.A(
        \PLUSE_0/bri_state_0/csse_2_0_a4_2_11 ), .B(
        \PLUSE_0/bri_state_0/N_183 ), .C(
        \PLUSE_0/bri_state_0/csse_2_0_1 ), .Y(
        \PLUSE_0/bri_state_0/cs_ns_e[3] ));
    DFN1E1 \top_code_0/cal_data[4]  (.D(\GPMI_0_dataout[4] ), .CLK(
        GLA_net_1), .E(\top_code_0/cal_data_1_sqmuxa ), .Q(
        \top_code_0_cal_data[4] ));
    NOR2B \state_1ms_0/timecount_RNO_6[9]  (.A(
        \state_1ms_0/PLUSETIME[9]_net_1 ), .B(
        \state_1ms_0/CS[5]_net_1 ), .Y(\state_1ms_0/PLUSETIME_m[9] ));
    DFN1E1 \scalestate_0/PLUSETIME180[1]  (.D(
        \top_code_0_scaledatain[1] ), .CLK(GLA_net_1), .E(
        \scalestate_0/PLUSETIME180_1_sqmuxa ), .Q(
        \scalestate_0/PLUSETIME180[1]_net_1 ));
    DFN1E1 \plusestate_0/PLUSETIME[8]  (.D(\top_code_0_plusedata[8] ), 
        .CLK(GLA_net_1), .E(\plusestate_0/DUMPTIME_0_sqmuxa_net_1 ), 
        .Q(\plusestate_0/PLUSETIME[8]_net_1 ));
    OR2B \DDS_0/dds_state_0/cs_RNI4SGF[6]  (.A(
        \DDS_0/dds_state_0/cs[6]_net_1 ), .B(\DDS_0/i[3] ), .Y(
        \DDS_0/dds_state_0/N_226 ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/un1_data_m59  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/data[2]_net_1 )
        , .B(\s_acq_change_0_s_stripnum[2] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/i2_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0/N_60_i ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[7]  (.D(
        \top_code_0_scaledatain[7] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[7]_net_1 ));
    NOR2B \scalestate_0/CS_RNI4P3V1[14]  (.A(\scalestate_0/N_1309 ), 
        .B(\scalestate_0/N_1196 ), .Y(\scalestate_0/N_1259 ));
    DFN1E1 \plusestate_0/timecount_1[14]  (.D(
        \plusestate_0/timecount_5[14] ), .CLK(GLA_net_1), .E(
        \plusestate_0/un1_sw_acq1_2_sqmuxa ), .Q(
        \plusestate_0_timecount[14] ));
    MX2 \top_code_0/inv_turn_RNO_0  (.A(top_code_0_inv_turn), .B(
        \xa_c[0] ), .S(\top_code_0/N_122 ), .Y(\top_code_0/N_802 ));
    DFN1 \state_1ms_0/timecount[13]  (.D(
        \state_1ms_0/timecount_RNO[13]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[13] ));
    XOR2 \DUMP_0/dump_coder_0/para3_RNIINFH[5]  (.A(
        \DUMP_0/dump_coder_0/para3[5]_net_1 ), .B(\DUMP_0/count_0[5] ), 
        .Y(\DUMP_0/dump_coder_0/un1_count_2_5[0] ));
    MX2 \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m92  (.A(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_91 ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_92 ), .S(
        \top_code_0_s_addchoice_0[1] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_93 ));
    DFN1 \state1ms_choice_0/dump_start  (.D(
        \state1ms_choice_0/dump_start_RNO_1 ), .CLK(GLA_net_1), .Q(
        state1ms_choice_0_dump_start));
    NOR2B \scalestate_0/necount_LE_NE_RNO  (.A(
        \scalestate_0/necount_LE_NE_1 ), .B(top_code_0_scale_rst_4), 
        .Y(\scalestate_0/necount_LE_NE_RNO_net_1 ));
    DFN1 \scalestate_0/strippluse[1]  (.D(
        \scalestate_0/strippluse_RNO[1]_net_1 ), .CLK(GLA_net_1), .Q(
        \scalestate_0_strippluse[1] ));
    NOR3C \scalestate_0/timecount_ret_28_RNO_7  (.A(
        top_code_0_scale_rst_0), .B(
        \scalestate_0/timecount_16_sqmuxa_1 ), .C(
        \scalestate_0/CUTTIME180_Tini[1]_net_1 ), .Y(
        \scalestate_0/CUTTIME180_Tini_m[1] ));
    AX1C \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_RNO[10]  (
        .A(\Signal_Noise_Acq_0/noise_acq_0/addr[9] ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_c8 ), .C(
        \Signal_Noise_Acq_0/noise_acq_0/addr[10] ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/noise_addr_1/addr_n10 ));
    NOR3C \sd_acq_top_0/sd_sacq_coder_0/i_RNO[6]  (.A(
        \sd_acq_top_0/sd_sacq_coder_0/i_reg18_NE[0] ), .B(
        \sd_acq_top_0/sd_sacq_coder_0/un1_count_4_NE[0] ), .C(
        \sd_acq_top_0/sd_sacq_coder_0/i_0_0[6] ), .Y(
        \sd_acq_top_0/sd_sacq_coder_0/i_RNO_0[6]_net_1 ));
    DFN1C0 \Signal_Noise_Acq_0/signal_acq_0/add_reg_5/addresult[3]  (
        .D(\Signal_Noise_Acq_0/signal_acq_0/add_reg_5/N_66_i ), .CLK(
        \Signal_Noise_Acq_0/signal_acq_0/signalclkctrl_0_clk_add ), 
        .CLR(s_acq_change_0_s_rst), .Q(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[3] ));
    DFN1C0 \PLUSE_0/bri_timer_0/count[5]/U1  (.D(
        \PLUSE_0/bri_timer_0/count[5]/Y ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .Q(\PLUSE_0/count_2[5] ));
    DFN1 \state_1ms_0/timecount[8]  (.D(
        \state_1ms_0/timecount_RNO[8]_net_1 ), .CLK(GLA_net_1), .Q(
        \state_1ms_0_timecount[8] ));
    DFN1E1 \top_code_0/state_1ms_data[14]  (.D(\GPMI_0_dataout[14] ), 
        .CLK(GLA_net_1), .E(\top_code_0/state_1ms_data_1_sqmuxa ), .Q(
        \top_code_0_state_1ms_data[14] ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_3[12]  (.A(
        \state_1ms_0_timecount[12] ), .B(
        \timer_top_0/state_switch_0/N_289 ), .Y(
        \timer_top_0/state_switch_0/N_257 ));
    MX2 \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_155  (.A(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR8_0_net ), .B(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/QX_TEMPR9_0_net ), .S(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/BUFF_11_Y ), .Y(
        \Signal_Noise_Acq_0/noise_acq_0/RAM_0/MX2_155_Y ));
    NOR3B \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/m213  (.A(
        \top_code_0_s_addchoice_3[0] ), .B(
        \Signal_Noise_Acq_0/signal_acq_0/addresult_1[9] ), .C(
        \top_code_0_s_addchoice_2[4] ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/rdata_choice_0/N_214 ));
    DFN1E1 \top_code_0/pd_pluse_data[4]  (.D(\GPMI_0_dataout_0[4] ), 
        .CLK(GLA_net_1), .E(\top_code_0/pd_pluse_data_1_sqmuxa ), .Q(
        \top_code_0_pd_pluse_data[4] ));
    XNOR3 
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/un3_addresult_m65  
        (.A(
        \Signal_Noise_Acq_0/signal_acq_0/un1_ten_choice_one_0_1[3] ), 
        .B(\Signal_Noise_Acq_0/signal_acq_0/addresult_4[3] ), .C(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/i4_mux ), .Y(
        \Signal_Noise_Acq_0/signal_acq_0/add_reg_1/N_66_i ));
    NOR2B \s_acq_change_0/s_stripnum_RNO[6]  (.A(\s_acq_change_0/N_62 )
        , .B(net_27), .Y(\s_acq_change_0/s_stripnum_RNO[6]_net_1 ));
    DFN1E1 \ClockManagement_0/long_timer_0/count[7]  (.D(
        \ClockManagement_0/long_timer_0/count_n7 ), .CLK(GLA_net_1), 
        .E(\ClockManagement_0/long_timer_0/counte ), .Q(
        \ClockManagement_0/long_timer_0/count[7]_net_1 ));
    NOR2B \top_code_0/relay_close_RNO[7]  (.A(\top_code_0/N_826 ), .B(
        net_27), .Y(\top_code_0/relay_close_RNO[7]_net_1 ));
    MX2 \state_1ms_0/timecount_RNO_0[0]  (.A(
        \state_1ms_0/timecount_8[0] ), .B(\state_1ms_0_timecount[0] ), 
        .S(\state_1ms_0/CS[9]_net_1 ), .Y(\state_1ms_0/N_67 ));
    XA1B \DUMP_0/dump_state_0/cs_srsts_0_0_a2_1[6]  (.A(\DUMP_0/i[6] ), 
        .B(\DUMP_0/i[4] ), .C(\DUMP_0/i[8] ), .Y(
        \DUMP_0/dump_state_0/N_203 ));
    NOR2B \timer_top_0/state_switch_0/dataout_RNO_4[2]  (.A(
        \plusestate_0_timecount[2] ), .B(
        \timer_top_0/state_switch_0/N_297 ), .Y(
        \timer_top_0/state_switch_0/N_234 ));
    DFN1E1 \state_1ms_0/CUTTIME[11]  (.D(
        \top_code_0_state_1ms_data[11] ), .CLK(GLA_net_1), .E(
        \state_1ms_0/N_364 ), .Q(\state_1ms_0/CUTTIME[11]_net_1 ));
    DFN1E1 \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[4]  (.D(
        \top_code_0_sd_sacq_data[4] ), .CLK(GLA_net_1), .E(
        \sd_acq_top_0/sd_sacq_coder_0/N_366 ), .Q(
        \sd_acq_top_0/sd_sacq_coder_0/sd_sacq_data5[4]_net_1 ));
    DFN1E1 \scalestate_0/CUTTIME180_TEL[14]  (.D(
        \top_code_0_scaledatain[14] ), .CLK(GLA_net_1), .E(
        \scalestate_0/N_1707 ), .Q(
        \scalestate_0/CUTTIME180_TEL[14]_net_1 ));
    DFN1E0 \DUMP_0/dump_coder_0/para5[9]  (.D(
        \DUMP_0/dump_coder_0/para5_4[9] ), .CLK(GLA_net_1), .E(
        \DUMP_0/dump_coder_0/un1_para114_2_net_1 ), .Q(
        \DUMP_0/dump_coder_0/para5[9]_net_1 ));
    DFN1E1 \DDS_0/dds_state_0/para_reg[5]  (.D(
        \top_code_0_dds_configdata[4] ), .CLK(GLA_net_1), .E(
        \DDS_0/dds_state_0/N_538_0 ), .Q(
        \DDS_0/dds_state_0/para_reg[5]_net_1 ));
    NOR2A \DUMP_0/dump_coder_0/para4_4[5]  (.A(
        \top_code_0_dumpdata_0[5] ), .B(\top_code_0_dump_cho_0[2] ), 
        .Y(\DUMP_0/dump_coder_0/para4_4[5]_net_1 ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
