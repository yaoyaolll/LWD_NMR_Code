`timescale 1 ns/100 ps
// Version: 9.1 9.1.0.18


module signal_acq(
       s_reset,
       signal_load,
       clk_sys,
       Signal_acq_clk,
       clk_dds,
       s_acq_en,
       acqnum,
       stripnum,
       s_periodnum,
       signal_data,
       s_addchoice,
       s_ADC
    );
input  s_reset;
input  signal_load;
input  clk_sys;
output Signal_acq_clk;
input  clk_dds;
input  s_acq_en;
input  [15:0] acqnum;
input  [11:0] stripnum;
input  [3:0] s_periodnum;
output [15:0] signal_data;
input  [4:0] s_addchoice;
input  [11:0] s_ADC;

    wire \add_reg_0_addresult_[19] , \add_reg_0_addresult_[18] , 
        \add_reg_0_addresult_[17] , \add_reg_0_addresult_[16] , 
        \add_reg_0_addresult_[15] , \add_reg_0_addresult_[14] , 
        \add_reg_0_addresult_[13] , \add_reg_0_addresult_[12] , 
        \add_reg_0_addresult_[11] , \add_reg_0_addresult_[10] , 
        \add_reg_0_addresult_[9] , \add_reg_0_addresult_[8] , 
        \add_reg_0_addresult_[7] , \add_reg_0_addresult_[6] , 
        \add_reg_0_addresult_[5] , \add_reg_0_addresult_[4] , 
        \add_reg_0_addresult_[3] , \add_reg_0_addresult_[2] , 
        \add_reg_0_addresult_[1] , \add_reg_0_addresult_[0] , 
        \add_reg_1_addresult_[19] , \add_reg_1_addresult_[18] , 
        \add_reg_1_addresult_[17] , \add_reg_1_addresult_[16] , 
        \add_reg_1_addresult_[15] , \add_reg_1_addresult_[14] , 
        \add_reg_1_addresult_[13] , \add_reg_1_addresult_[12] , 
        \add_reg_1_addresult_[11] , \add_reg_1_addresult_[10] , 
        \add_reg_1_addresult_[9] , \add_reg_1_addresult_[8] , 
        \add_reg_1_addresult_[7] , \add_reg_1_addresult_[6] , 
        \add_reg_1_addresult_[5] , \add_reg_1_addresult_[4] , 
        \add_reg_1_addresult_[3] , \add_reg_1_addresult_[2] , 
        \add_reg_1_addresult_[1] , \add_reg_1_addresult_[0] , 
        \add_reg_2_addresult_[19] , \add_reg_2_addresult_[18] , 
        \add_reg_2_addresult_[17] , \add_reg_2_addresult_[16] , 
        \add_reg_2_addresult_[15] , \add_reg_2_addresult_[14] , 
        \add_reg_2_addresult_[13] , \add_reg_2_addresult_[12] , 
        \add_reg_2_addresult_[11] , \add_reg_2_addresult_[10] , 
        \add_reg_2_addresult_[9] , \add_reg_2_addresult_[8] , 
        \add_reg_2_addresult_[7] , \add_reg_2_addresult_[6] , 
        \add_reg_2_addresult_[5] , \add_reg_2_addresult_[4] , 
        \add_reg_2_addresult_[3] , \add_reg_2_addresult_[2] , 
        \add_reg_2_addresult_[1] , \add_reg_2_addresult_[0] , 
        \add_reg_3_addresult_[19] , \add_reg_3_addresult_[18] , 
        \add_reg_3_addresult_[17] , \add_reg_3_addresult_[16] , 
        \add_reg_3_addresult_[15] , \add_reg_3_addresult_[14] , 
        \add_reg_3_addresult_[13] , \add_reg_3_addresult_[12] , 
        \add_reg_3_addresult_[11] , \add_reg_3_addresult_[10] , 
        \add_reg_3_addresult_[9] , \add_reg_3_addresult_[8] , 
        \add_reg_3_addresult_[7] , \add_reg_3_addresult_[6] , 
        \add_reg_3_addresult_[5] , \add_reg_3_addresult_[4] , 
        \add_reg_3_addresult_[3] , \add_reg_3_addresult_[2] , 
        \add_reg_3_addresult_[1] , \add_reg_3_addresult_[0] , 
        \add_reg_4_addresult_[19] , \add_reg_4_addresult_[18] , 
        \add_reg_4_addresult_[17] , \add_reg_4_addresult_[16] , 
        \add_reg_4_addresult_[15] , \add_reg_4_addresult_[14] , 
        \add_reg_4_addresult_[13] , \add_reg_4_addresult_[12] , 
        \add_reg_4_addresult_[11] , \add_reg_4_addresult_[10] , 
        \add_reg_4_addresult_[9] , \add_reg_4_addresult_[8] , 
        \add_reg_4_addresult_[7] , \add_reg_4_addresult_[6] , 
        \add_reg_4_addresult_[5] , \add_reg_4_addresult_[4] , 
        \add_reg_4_addresult_[3] , \add_reg_4_addresult_[2] , 
        \add_reg_4_addresult_[1] , \add_reg_4_addresult_[0] , 
        \add_reg_5_addresult_[19] , \add_reg_5_addresult_[18] , 
        \add_reg_5_addresult_[17] , \add_reg_5_addresult_[16] , 
        \add_reg_5_addresult_[15] , \add_reg_5_addresult_[14] , 
        \add_reg_5_addresult_[13] , \add_reg_5_addresult_[12] , 
        \add_reg_5_addresult_[11] , \add_reg_5_addresult_[10] , 
        \add_reg_5_addresult_[9] , \add_reg_5_addresult_[8] , 
        \add_reg_5_addresult_[7] , \add_reg_5_addresult_[6] , 
        \add_reg_5_addresult_[5] , \add_reg_5_addresult_[4] , 
        \add_reg_5_addresult_[3] , \add_reg_5_addresult_[2] , 
        \add_reg_5_addresult_[1] , \add_reg_5_addresult_[0] , 
        \add_reg_6_addresult_[19] , \add_reg_6_addresult_[18] , 
        \add_reg_6_addresult_[17] , \add_reg_6_addresult_[16] , 
        \add_reg_6_addresult_[15] , \add_reg_6_addresult_[14] , 
        \add_reg_6_addresult_[13] , \add_reg_6_addresult_[12] , 
        \add_reg_6_addresult_[11] , \add_reg_6_addresult_[10] , 
        \add_reg_6_addresult_[9] , \add_reg_6_addresult_[8] , 
        \add_reg_6_addresult_[7] , \add_reg_6_addresult_[6] , 
        \add_reg_6_addresult_[5] , \add_reg_6_addresult_[4] , 
        \add_reg_6_addresult_[3] , \add_reg_6_addresult_[2] , 
        \add_reg_6_addresult_[1] , \add_reg_6_addresult_[0] , 
        \add_reg_7_addresult_[19] , \add_reg_7_addresult_[18] , 
        \add_reg_7_addresult_[17] , \add_reg_7_addresult_[16] , 
        \add_reg_7_addresult_[15] , \add_reg_7_addresult_[14] , 
        \add_reg_7_addresult_[13] , \add_reg_7_addresult_[12] , 
        \add_reg_7_addresult_[11] , \add_reg_7_addresult_[10] , 
        \add_reg_7_addresult_[9] , \add_reg_7_addresult_[8] , 
        \add_reg_7_addresult_[7] , \add_reg_7_addresult_[6] , 
        \add_reg_7_addresult_[5] , \add_reg_7_addresult_[4] , 
        \add_reg_7_addresult_[3] , \add_reg_7_addresult_[2] , 
        \add_reg_7_addresult_[1] , \add_reg_7_addresult_[0] , 
        \ctrl_addr_0_addrout_[3] , \ctrl_addr_0_addrout_[2] , 
        \ctrl_addr_0_addrout_[1] , \ctrl_addr_0_addrout_[0] , 
        signalclkctrl_0_clk_add, signalclkctrl_0_entop, 
        s_clk_div4_0_clkout, \ten_choice_one_0_dataeight_[11] , 
        \ten_choice_one_0_dataeight_[10] , 
        \ten_choice_one_0_dataeight_[9] , 
        \ten_choice_one_0_dataeight_[8] , 
        \ten_choice_one_0_dataeight_[7] , 
        \ten_choice_one_0_dataeight_[6] , 
        \ten_choice_one_0_dataeight_[5] , 
        \ten_choice_one_0_dataeight_[4] , 
        \ten_choice_one_0_dataeight_[3] , 
        \ten_choice_one_0_dataeight_[2] , 
        \ten_choice_one_0_dataeight_[1] , 
        \ten_choice_one_0_dataeight_[0] , 
        \ten_choice_one_0_datafive_[11] , 
        \ten_choice_one_0_datafive_[10] , 
        \ten_choice_one_0_datafive_[9] , 
        \ten_choice_one_0_datafive_[8] , 
        \ten_choice_one_0_datafive_[7] , 
        \ten_choice_one_0_datafive_[6] , 
        \ten_choice_one_0_datafive_[5] , 
        \ten_choice_one_0_datafive_[4] , 
        \ten_choice_one_0_datafive_[3] , 
        \ten_choice_one_0_datafive_[2] , 
        \ten_choice_one_0_datafive_[1] , 
        \ten_choice_one_0_datafive_[0] , 
        \ten_choice_one_0_datafour_[11] , 
        \ten_choice_one_0_datafour_[10] , 
        \ten_choice_one_0_datafour_[9] , 
        \ten_choice_one_0_datafour_[8] , 
        \ten_choice_one_0_datafour_[7] , 
        \ten_choice_one_0_datafour_[6] , 
        \ten_choice_one_0_datafour_[5] , 
        \ten_choice_one_0_datafour_[4] , 
        \ten_choice_one_0_datafour_[3] , 
        \ten_choice_one_0_datafour_[2] , 
        \ten_choice_one_0_datafour_[1] , 
        \ten_choice_one_0_datafour_[0] , 
        \ten_choice_one_0_dataone_[11] , 
        \ten_choice_one_0_dataone_[10] , 
        \ten_choice_one_0_dataone_[9] , \ten_choice_one_0_dataone_[8] , 
        \ten_choice_one_0_dataone_[7] , \ten_choice_one_0_dataone_[6] , 
        \ten_choice_one_0_dataone_[5] , \ten_choice_one_0_dataone_[4] , 
        \ten_choice_one_0_dataone_[3] , \ten_choice_one_0_dataone_[2] , 
        \ten_choice_one_0_dataone_[1] , \ten_choice_one_0_dataone_[0] , 
        \ten_choice_one_0_dataseven_[11] , 
        \ten_choice_one_0_dataseven_[10] , 
        \ten_choice_one_0_dataseven_[9] , 
        \ten_choice_one_0_dataseven_[8] , 
        \ten_choice_one_0_dataseven_[7] , 
        \ten_choice_one_0_dataseven_[6] , 
        \ten_choice_one_0_dataseven_[5] , 
        \ten_choice_one_0_dataseven_[4] , 
        \ten_choice_one_0_dataseven_[3] , 
        \ten_choice_one_0_dataseven_[2] , 
        \ten_choice_one_0_dataseven_[1] , 
        \ten_choice_one_0_dataseven_[0] , 
        \ten_choice_one_0_datasix_[11] , 
        \ten_choice_one_0_datasix_[10] , 
        \ten_choice_one_0_datasix_[9] , \ten_choice_one_0_datasix_[8] , 
        \ten_choice_one_0_datasix_[7] , \ten_choice_one_0_datasix_[6] , 
        \ten_choice_one_0_datasix_[5] , \ten_choice_one_0_datasix_[4] , 
        \ten_choice_one_0_datasix_[3] , \ten_choice_one_0_datasix_[2] , 
        \ten_choice_one_0_datasix_[1] , \ten_choice_one_0_datasix_[0] , 
        \ten_choice_one_0_datathree_[11] , 
        \ten_choice_one_0_datathree_[10] , 
        \ten_choice_one_0_datathree_[9] , 
        \ten_choice_one_0_datathree_[8] , 
        \ten_choice_one_0_datathree_[7] , 
        \ten_choice_one_0_datathree_[6] , 
        \ten_choice_one_0_datathree_[5] , 
        \ten_choice_one_0_datathree_[4] , 
        \ten_choice_one_0_datathree_[3] , 
        \ten_choice_one_0_datathree_[2] , 
        \ten_choice_one_0_datathree_[1] , 
        \ten_choice_one_0_datathree_[0] , 
        \ten_choice_one_0_datatwo_[11] , 
        \ten_choice_one_0_datatwo_[10] , 
        \ten_choice_one_0_datatwo_[9] , \ten_choice_one_0_datatwo_[8] , 
        \ten_choice_one_0_datatwo_[7] , \ten_choice_one_0_datatwo_[6] , 
        \ten_choice_one_0_datatwo_[5] , \ten_choice_one_0_datatwo_[4] , 
        \ten_choice_one_0_datatwo_[3] , \ten_choice_one_0_datatwo_[2] , 
        \ten_choice_one_0_datatwo_[1] , \ten_choice_one_0_datatwo_[0] , 
        GND_net, VCC_net;
    
    add_reg add_reg_2 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_datathree_[11] , 
        \ten_choice_one_0_datathree_[10] , 
        \ten_choice_one_0_datathree_[9] , 
        \ten_choice_one_0_datathree_[8] , 
        \ten_choice_one_0_datathree_[7] , 
        \ten_choice_one_0_datathree_[6] , 
        \ten_choice_one_0_datathree_[5] , 
        \ten_choice_one_0_datathree_[4] , 
        \ten_choice_one_0_datathree_[3] , 
        \ten_choice_one_0_datathree_[2] , 
        \ten_choice_one_0_datathree_[1] , 
        \ten_choice_one_0_datathree_[0] }), .addresult({
        \add_reg_2_addresult_[19] , \add_reg_2_addresult_[18] , 
        \add_reg_2_addresult_[17] , \add_reg_2_addresult_[16] , 
        \add_reg_2_addresult_[15] , \add_reg_2_addresult_[14] , 
        \add_reg_2_addresult_[13] , \add_reg_2_addresult_[12] , 
        \add_reg_2_addresult_[11] , \add_reg_2_addresult_[10] , 
        \add_reg_2_addresult_[9] , \add_reg_2_addresult_[8] , 
        \add_reg_2_addresult_[7] , \add_reg_2_addresult_[6] , 
        \add_reg_2_addresult_[5] , \add_reg_2_addresult_[4] , 
        \add_reg_2_addresult_[3] , \add_reg_2_addresult_[2] , 
        \add_reg_2_addresult_[1] , \add_reg_2_addresult_[0] }));
    s_clk_div4 s_clk_div4_0 (.rst_n(s_reset), .entop(
        signalclkctrl_0_entop), .s_acq_en(s_acq_en), .clk_dds(clk_dds), 
        .clkout(s_clk_div4_0_clkout));
    signalclkctrl signalclkctrl_0 (.rst_n(s_reset), .clk_sys(clk_sys), 
        .load(signal_load), .entop(signalclkctrl_0_entop), .clk_add(
        signalclkctrl_0_clk_add), .clk_acq(Signal_acq_clk), .clkin(
        s_clk_div4_0_clkout), .acqnum({acqnum[15], acqnum[14], 
        acqnum[13], acqnum[12], acqnum[11], acqnum[10], acqnum[9], 
        acqnum[8], acqnum[7], acqnum[6], acqnum[5], acqnum[4], 
        acqnum[3], acqnum[2], acqnum[1], acqnum[0]}), .stripnum({
        stripnum[11], stripnum[10], stripnum[9], stripnum[8], 
        stripnum[7], stripnum[6], stripnum[5], stripnum[4], 
        stripnum[3], stripnum[2], stripnum[1], stripnum[0]}), 
        .periodnum({s_periodnum[3], s_periodnum[2], s_periodnum[1], 
        s_periodnum[0]}));
    rdata_choice rdata_choice_0 (.dataone({\add_reg_0_addresult_[19] , 
        \add_reg_0_addresult_[18] , \add_reg_0_addresult_[17] , 
        \add_reg_0_addresult_[16] , \add_reg_0_addresult_[15] , 
        \add_reg_0_addresult_[14] , \add_reg_0_addresult_[13] , 
        \add_reg_0_addresult_[12] , \add_reg_0_addresult_[11] , 
        \add_reg_0_addresult_[10] , \add_reg_0_addresult_[9] , 
        \add_reg_0_addresult_[8] , \add_reg_0_addresult_[7] , 
        \add_reg_0_addresult_[6] , \add_reg_0_addresult_[5] , 
        \add_reg_0_addresult_[4] , \add_reg_0_addresult_[3] , 
        \add_reg_0_addresult_[2] , \add_reg_0_addresult_[1] , 
        \add_reg_0_addresult_[0] }), .datatwo({
        \add_reg_1_addresult_[19] , \add_reg_1_addresult_[18] , 
        \add_reg_1_addresult_[17] , \add_reg_1_addresult_[16] , 
        \add_reg_1_addresult_[15] , \add_reg_1_addresult_[14] , 
        \add_reg_1_addresult_[13] , \add_reg_1_addresult_[12] , 
        \add_reg_1_addresult_[11] , \add_reg_1_addresult_[10] , 
        \add_reg_1_addresult_[9] , \add_reg_1_addresult_[8] , 
        \add_reg_1_addresult_[7] , \add_reg_1_addresult_[6] , 
        \add_reg_1_addresult_[5] , \add_reg_1_addresult_[4] , 
        \add_reg_1_addresult_[3] , \add_reg_1_addresult_[2] , 
        \add_reg_1_addresult_[1] , \add_reg_1_addresult_[0] }), 
        .datathree({\add_reg_2_addresult_[19] , 
        \add_reg_2_addresult_[18] , \add_reg_2_addresult_[17] , 
        \add_reg_2_addresult_[16] , \add_reg_2_addresult_[15] , 
        \add_reg_2_addresult_[14] , \add_reg_2_addresult_[13] , 
        \add_reg_2_addresult_[12] , \add_reg_2_addresult_[11] , 
        \add_reg_2_addresult_[10] , \add_reg_2_addresult_[9] , 
        \add_reg_2_addresult_[8] , \add_reg_2_addresult_[7] , 
        \add_reg_2_addresult_[6] , \add_reg_2_addresult_[5] , 
        \add_reg_2_addresult_[4] , \add_reg_2_addresult_[3] , 
        \add_reg_2_addresult_[2] , \add_reg_2_addresult_[1] , 
        \add_reg_2_addresult_[0] }), .datafour({
        \add_reg_3_addresult_[19] , \add_reg_3_addresult_[18] , 
        \add_reg_3_addresult_[17] , \add_reg_3_addresult_[16] , 
        \add_reg_3_addresult_[15] , \add_reg_3_addresult_[14] , 
        \add_reg_3_addresult_[13] , \add_reg_3_addresult_[12] , 
        \add_reg_3_addresult_[11] , \add_reg_3_addresult_[10] , 
        \add_reg_3_addresult_[9] , \add_reg_3_addresult_[8] , 
        \add_reg_3_addresult_[7] , \add_reg_3_addresult_[6] , 
        \add_reg_3_addresult_[5] , \add_reg_3_addresult_[4] , 
        \add_reg_3_addresult_[3] , \add_reg_3_addresult_[2] , 
        \add_reg_3_addresult_[1] , \add_reg_3_addresult_[0] }), 
        .datafive({\add_reg_4_addresult_[19] , 
        \add_reg_4_addresult_[18] , \add_reg_4_addresult_[17] , 
        \add_reg_4_addresult_[16] , \add_reg_4_addresult_[15] , 
        \add_reg_4_addresult_[14] , \add_reg_4_addresult_[13] , 
        \add_reg_4_addresult_[12] , \add_reg_4_addresult_[11] , 
        \add_reg_4_addresult_[10] , \add_reg_4_addresult_[9] , 
        \add_reg_4_addresult_[8] , \add_reg_4_addresult_[7] , 
        \add_reg_4_addresult_[6] , \add_reg_4_addresult_[5] , 
        \add_reg_4_addresult_[4] , \add_reg_4_addresult_[3] , 
        \add_reg_4_addresult_[2] , \add_reg_4_addresult_[1] , 
        \add_reg_4_addresult_[0] }), .datasix({
        \add_reg_5_addresult_[19] , \add_reg_5_addresult_[18] , 
        \add_reg_5_addresult_[17] , \add_reg_5_addresult_[16] , 
        \add_reg_5_addresult_[15] , \add_reg_5_addresult_[14] , 
        \add_reg_5_addresult_[13] , \add_reg_5_addresult_[12] , 
        \add_reg_5_addresult_[11] , \add_reg_5_addresult_[10] , 
        \add_reg_5_addresult_[9] , \add_reg_5_addresult_[8] , 
        \add_reg_5_addresult_[7] , \add_reg_5_addresult_[6] , 
        \add_reg_5_addresult_[5] , \add_reg_5_addresult_[4] , 
        \add_reg_5_addresult_[3] , \add_reg_5_addresult_[2] , 
        \add_reg_5_addresult_[1] , \add_reg_5_addresult_[0] }), 
        .dataseven({\add_reg_6_addresult_[19] , 
        \add_reg_6_addresult_[18] , \add_reg_6_addresult_[17] , 
        \add_reg_6_addresult_[16] , \add_reg_6_addresult_[15] , 
        \add_reg_6_addresult_[14] , \add_reg_6_addresult_[13] , 
        \add_reg_6_addresult_[12] , \add_reg_6_addresult_[11] , 
        \add_reg_6_addresult_[10] , \add_reg_6_addresult_[9] , 
        \add_reg_6_addresult_[8] , \add_reg_6_addresult_[7] , 
        \add_reg_6_addresult_[6] , \add_reg_6_addresult_[5] , 
        \add_reg_6_addresult_[4] , \add_reg_6_addresult_[3] , 
        \add_reg_6_addresult_[2] , \add_reg_6_addresult_[1] , 
        \add_reg_6_addresult_[0] }), .dataeight({
        \add_reg_7_addresult_[19] , \add_reg_7_addresult_[18] , 
        \add_reg_7_addresult_[17] , \add_reg_7_addresult_[16] , 
        \add_reg_7_addresult_[15] , \add_reg_7_addresult_[14] , 
        \add_reg_7_addresult_[13] , \add_reg_7_addresult_[12] , 
        \add_reg_7_addresult_[11] , \add_reg_7_addresult_[10] , 
        \add_reg_7_addresult_[9] , \add_reg_7_addresult_[8] , 
        \add_reg_7_addresult_[7] , \add_reg_7_addresult_[6] , 
        \add_reg_7_addresult_[5] , \add_reg_7_addresult_[4] , 
        \add_reg_7_addresult_[3] , \add_reg_7_addresult_[2] , 
        \add_reg_7_addresult_[1] , \add_reg_7_addresult_[0] }), 
        .dataout({signal_data[15], signal_data[14], signal_data[13], 
        signal_data[12], signal_data[11], signal_data[10], 
        signal_data[9], signal_data[8], signal_data[7], signal_data[6], 
        signal_data[5], signal_data[4], signal_data[3], signal_data[2], 
        signal_data[1], signal_data[0]}), .choice({s_addchoice[4], 
        s_addchoice[3], s_addchoice[2], s_addchoice[1], s_addchoice[0]})
        );
    GND GND (.Y(GND_net));
    add_reg add_reg_5 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_datasix_[11] , 
        \ten_choice_one_0_datasix_[10] , 
        \ten_choice_one_0_datasix_[9] , \ten_choice_one_0_datasix_[8] , 
        \ten_choice_one_0_datasix_[7] , \ten_choice_one_0_datasix_[6] , 
        \ten_choice_one_0_datasix_[5] , \ten_choice_one_0_datasix_[4] , 
        \ten_choice_one_0_datasix_[3] , \ten_choice_one_0_datasix_[2] , 
        \ten_choice_one_0_datasix_[1] , \ten_choice_one_0_datasix_[0] })
        , .addresult({\add_reg_5_addresult_[19] , 
        \add_reg_5_addresult_[18] , \add_reg_5_addresult_[17] , 
        \add_reg_5_addresult_[16] , \add_reg_5_addresult_[15] , 
        \add_reg_5_addresult_[14] , \add_reg_5_addresult_[13] , 
        \add_reg_5_addresult_[12] , \add_reg_5_addresult_[11] , 
        \add_reg_5_addresult_[10] , \add_reg_5_addresult_[9] , 
        \add_reg_5_addresult_[8] , \add_reg_5_addresult_[7] , 
        \add_reg_5_addresult_[6] , \add_reg_5_addresult_[5] , 
        \add_reg_5_addresult_[4] , \add_reg_5_addresult_[3] , 
        \add_reg_5_addresult_[2] , \add_reg_5_addresult_[1] , 
        \add_reg_5_addresult_[0] }));
    add_reg add_reg_3 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_datafour_[11] , 
        \ten_choice_one_0_datafour_[10] , 
        \ten_choice_one_0_datafour_[9] , 
        \ten_choice_one_0_datafour_[8] , 
        \ten_choice_one_0_datafour_[7] , 
        \ten_choice_one_0_datafour_[6] , 
        \ten_choice_one_0_datafour_[5] , 
        \ten_choice_one_0_datafour_[4] , 
        \ten_choice_one_0_datafour_[3] , 
        \ten_choice_one_0_datafour_[2] , 
        \ten_choice_one_0_datafour_[1] , 
        \ten_choice_one_0_datafour_[0] }), .addresult({
        \add_reg_3_addresult_[19] , \add_reg_3_addresult_[18] , 
        \add_reg_3_addresult_[17] , \add_reg_3_addresult_[16] , 
        \add_reg_3_addresult_[15] , \add_reg_3_addresult_[14] , 
        \add_reg_3_addresult_[13] , \add_reg_3_addresult_[12] , 
        \add_reg_3_addresult_[11] , \add_reg_3_addresult_[10] , 
        \add_reg_3_addresult_[9] , \add_reg_3_addresult_[8] , 
        \add_reg_3_addresult_[7] , \add_reg_3_addresult_[6] , 
        \add_reg_3_addresult_[5] , \add_reg_3_addresult_[4] , 
        \add_reg_3_addresult_[3] , \add_reg_3_addresult_[2] , 
        \add_reg_3_addresult_[1] , \add_reg_3_addresult_[0] }));
    add_reg add_reg_1 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_datatwo_[11] , 
        \ten_choice_one_0_datatwo_[10] , 
        \ten_choice_one_0_datatwo_[9] , \ten_choice_one_0_datatwo_[8] , 
        \ten_choice_one_0_datatwo_[7] , \ten_choice_one_0_datatwo_[6] , 
        \ten_choice_one_0_datatwo_[5] , \ten_choice_one_0_datatwo_[4] , 
        \ten_choice_one_0_datatwo_[3] , \ten_choice_one_0_datatwo_[2] , 
        \ten_choice_one_0_datatwo_[1] , \ten_choice_one_0_datatwo_[0] })
        , .addresult({\add_reg_1_addresult_[19] , 
        \add_reg_1_addresult_[18] , \add_reg_1_addresult_[17] , 
        \add_reg_1_addresult_[16] , \add_reg_1_addresult_[15] , 
        \add_reg_1_addresult_[14] , \add_reg_1_addresult_[13] , 
        \add_reg_1_addresult_[12] , \add_reg_1_addresult_[11] , 
        \add_reg_1_addresult_[10] , \add_reg_1_addresult_[9] , 
        \add_reg_1_addresult_[8] , \add_reg_1_addresult_[7] , 
        \add_reg_1_addresult_[6] , \add_reg_1_addresult_[5] , 
        \add_reg_1_addresult_[4] , \add_reg_1_addresult_[3] , 
        \add_reg_1_addresult_[2] , \add_reg_1_addresult_[1] , 
        \add_reg_1_addresult_[0] }));
    add_reg add_reg_0 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_dataone_[11] , 
        \ten_choice_one_0_dataone_[10] , 
        \ten_choice_one_0_dataone_[9] , \ten_choice_one_0_dataone_[8] , 
        \ten_choice_one_0_dataone_[7] , \ten_choice_one_0_dataone_[6] , 
        \ten_choice_one_0_dataone_[5] , \ten_choice_one_0_dataone_[4] , 
        \ten_choice_one_0_dataone_[3] , \ten_choice_one_0_dataone_[2] , 
        \ten_choice_one_0_dataone_[1] , \ten_choice_one_0_dataone_[0] })
        , .addresult({\add_reg_0_addresult_[19] , 
        \add_reg_0_addresult_[18] , \add_reg_0_addresult_[17] , 
        \add_reg_0_addresult_[16] , \add_reg_0_addresult_[15] , 
        \add_reg_0_addresult_[14] , \add_reg_0_addresult_[13] , 
        \add_reg_0_addresult_[12] , \add_reg_0_addresult_[11] , 
        \add_reg_0_addresult_[10] , \add_reg_0_addresult_[9] , 
        \add_reg_0_addresult_[8] , \add_reg_0_addresult_[7] , 
        \add_reg_0_addresult_[6] , \add_reg_0_addresult_[5] , 
        \add_reg_0_addresult_[4] , \add_reg_0_addresult_[3] , 
        \add_reg_0_addresult_[2] , \add_reg_0_addresult_[1] , 
        \add_reg_0_addresult_[0] }));
    VCC VCC (.Y(VCC_net));
    ctrl_addr ctrl_addr_0 (.rst_n(s_reset), .clk_sys(clk_sys), .clk(
        signalclkctrl_0_clk_add), .load(signal_load), .addrout({
        \ctrl_addr_0_addrout_[3] , \ctrl_addr_0_addrout_[2] , 
        \ctrl_addr_0_addrout_[1] , \ctrl_addr_0_addrout_[0] }), 
        .datain({s_periodnum[3], s_periodnum[2], s_periodnum[1], 
        s_periodnum[0]}));
    add_reg add_reg_7 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_dataeight_[11] , 
        \ten_choice_one_0_dataeight_[10] , 
        \ten_choice_one_0_dataeight_[9] , 
        \ten_choice_one_0_dataeight_[8] , 
        \ten_choice_one_0_dataeight_[7] , 
        \ten_choice_one_0_dataeight_[6] , 
        \ten_choice_one_0_dataeight_[5] , 
        \ten_choice_one_0_dataeight_[4] , 
        \ten_choice_one_0_dataeight_[3] , 
        \ten_choice_one_0_dataeight_[2] , 
        \ten_choice_one_0_dataeight_[1] , 
        \ten_choice_one_0_dataeight_[0] }), .addresult({
        \add_reg_7_addresult_[19] , \add_reg_7_addresult_[18] , 
        \add_reg_7_addresult_[17] , \add_reg_7_addresult_[16] , 
        \add_reg_7_addresult_[15] , \add_reg_7_addresult_[14] , 
        \add_reg_7_addresult_[13] , \add_reg_7_addresult_[12] , 
        \add_reg_7_addresult_[11] , \add_reg_7_addresult_[10] , 
        \add_reg_7_addresult_[9] , \add_reg_7_addresult_[8] , 
        \add_reg_7_addresult_[7] , \add_reg_7_addresult_[6] , 
        \add_reg_7_addresult_[5] , \add_reg_7_addresult_[4] , 
        \add_reg_7_addresult_[3] , \add_reg_7_addresult_[2] , 
        \add_reg_7_addresult_[1] , \add_reg_7_addresult_[0] }));
    add_reg add_reg_6 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_dataseven_[11] , 
        \ten_choice_one_0_dataseven_[10] , 
        \ten_choice_one_0_dataseven_[9] , 
        \ten_choice_one_0_dataseven_[8] , 
        \ten_choice_one_0_dataseven_[7] , 
        \ten_choice_one_0_dataseven_[6] , 
        \ten_choice_one_0_dataseven_[5] , 
        \ten_choice_one_0_dataseven_[4] , 
        \ten_choice_one_0_dataseven_[3] , 
        \ten_choice_one_0_dataseven_[2] , 
        \ten_choice_one_0_dataseven_[1] , 
        \ten_choice_one_0_dataseven_[0] }), .addresult({
        \add_reg_6_addresult_[19] , \add_reg_6_addresult_[18] , 
        \add_reg_6_addresult_[17] , \add_reg_6_addresult_[16] , 
        \add_reg_6_addresult_[15] , \add_reg_6_addresult_[14] , 
        \add_reg_6_addresult_[13] , \add_reg_6_addresult_[12] , 
        \add_reg_6_addresult_[11] , \add_reg_6_addresult_[10] , 
        \add_reg_6_addresult_[9] , \add_reg_6_addresult_[8] , 
        \add_reg_6_addresult_[7] , \add_reg_6_addresult_[6] , 
        \add_reg_6_addresult_[5] , \add_reg_6_addresult_[4] , 
        \add_reg_6_addresult_[3] , \add_reg_6_addresult_[2] , 
        \add_reg_6_addresult_[1] , \add_reg_6_addresult_[0] }));
    add_reg add_reg_4 (.clk(signalclkctrl_0_clk_add), .rst_n(s_reset), 
        .addin({\ten_choice_one_0_datafive_[11] , 
        \ten_choice_one_0_datafive_[10] , 
        \ten_choice_one_0_datafive_[9] , 
        \ten_choice_one_0_datafive_[8] , 
        \ten_choice_one_0_datafive_[7] , 
        \ten_choice_one_0_datafive_[6] , 
        \ten_choice_one_0_datafive_[5] , 
        \ten_choice_one_0_datafive_[4] , 
        \ten_choice_one_0_datafive_[3] , 
        \ten_choice_one_0_datafive_[2] , 
        \ten_choice_one_0_datafive_[1] , 
        \ten_choice_one_0_datafive_[0] }), .addresult({
        \add_reg_4_addresult_[19] , \add_reg_4_addresult_[18] , 
        \add_reg_4_addresult_[17] , \add_reg_4_addresult_[16] , 
        \add_reg_4_addresult_[15] , \add_reg_4_addresult_[14] , 
        \add_reg_4_addresult_[13] , \add_reg_4_addresult_[12] , 
        \add_reg_4_addresult_[11] , \add_reg_4_addresult_[10] , 
        \add_reg_4_addresult_[9] , \add_reg_4_addresult_[8] , 
        \add_reg_4_addresult_[7] , \add_reg_4_addresult_[6] , 
        \add_reg_4_addresult_[5] , \add_reg_4_addresult_[4] , 
        \add_reg_4_addresult_[3] , \add_reg_4_addresult_[2] , 
        \add_reg_4_addresult_[1] , \add_reg_4_addresult_[0] }));
    ten_choice_one ten_choice_one_0 (.choice({
        \ctrl_addr_0_addrout_[3] , \ctrl_addr_0_addrout_[2] , 
        \ctrl_addr_0_addrout_[1] , \ctrl_addr_0_addrout_[0] }), 
        .dataone({\ten_choice_one_0_dataone_[11] , 
        \ten_choice_one_0_dataone_[10] , 
        \ten_choice_one_0_dataone_[9] , \ten_choice_one_0_dataone_[8] , 
        \ten_choice_one_0_dataone_[7] , \ten_choice_one_0_dataone_[6] , 
        \ten_choice_one_0_dataone_[5] , \ten_choice_one_0_dataone_[4] , 
        \ten_choice_one_0_dataone_[3] , \ten_choice_one_0_dataone_[2] , 
        \ten_choice_one_0_dataone_[1] , \ten_choice_one_0_dataone_[0] })
        , .datatwo({\ten_choice_one_0_datatwo_[11] , 
        \ten_choice_one_0_datatwo_[10] , 
        \ten_choice_one_0_datatwo_[9] , \ten_choice_one_0_datatwo_[8] , 
        \ten_choice_one_0_datatwo_[7] , \ten_choice_one_0_datatwo_[6] , 
        \ten_choice_one_0_datatwo_[5] , \ten_choice_one_0_datatwo_[4] , 
        \ten_choice_one_0_datatwo_[3] , \ten_choice_one_0_datatwo_[2] , 
        \ten_choice_one_0_datatwo_[1] , \ten_choice_one_0_datatwo_[0] })
        , .datathree({\ten_choice_one_0_datathree_[11] , 
        \ten_choice_one_0_datathree_[10] , 
        \ten_choice_one_0_datathree_[9] , 
        \ten_choice_one_0_datathree_[8] , 
        \ten_choice_one_0_datathree_[7] , 
        \ten_choice_one_0_datathree_[6] , 
        \ten_choice_one_0_datathree_[5] , 
        \ten_choice_one_0_datathree_[4] , 
        \ten_choice_one_0_datathree_[3] , 
        \ten_choice_one_0_datathree_[2] , 
        \ten_choice_one_0_datathree_[1] , 
        \ten_choice_one_0_datathree_[0] }), .datafour({
        \ten_choice_one_0_datafour_[11] , 
        \ten_choice_one_0_datafour_[10] , 
        \ten_choice_one_0_datafour_[9] , 
        \ten_choice_one_0_datafour_[8] , 
        \ten_choice_one_0_datafour_[7] , 
        \ten_choice_one_0_datafour_[6] , 
        \ten_choice_one_0_datafour_[5] , 
        \ten_choice_one_0_datafour_[4] , 
        \ten_choice_one_0_datafour_[3] , 
        \ten_choice_one_0_datafour_[2] , 
        \ten_choice_one_0_datafour_[1] , 
        \ten_choice_one_0_datafour_[0] }), .datafive({
        \ten_choice_one_0_datafive_[11] , 
        \ten_choice_one_0_datafive_[10] , 
        \ten_choice_one_0_datafive_[9] , 
        \ten_choice_one_0_datafive_[8] , 
        \ten_choice_one_0_datafive_[7] , 
        \ten_choice_one_0_datafive_[6] , 
        \ten_choice_one_0_datafive_[5] , 
        \ten_choice_one_0_datafive_[4] , 
        \ten_choice_one_0_datafive_[3] , 
        \ten_choice_one_0_datafive_[2] , 
        \ten_choice_one_0_datafive_[1] , 
        \ten_choice_one_0_datafive_[0] }), .datasix({
        \ten_choice_one_0_datasix_[11] , 
        \ten_choice_one_0_datasix_[10] , 
        \ten_choice_one_0_datasix_[9] , \ten_choice_one_0_datasix_[8] , 
        \ten_choice_one_0_datasix_[7] , \ten_choice_one_0_datasix_[6] , 
        \ten_choice_one_0_datasix_[5] , \ten_choice_one_0_datasix_[4] , 
        \ten_choice_one_0_datasix_[3] , \ten_choice_one_0_datasix_[2] , 
        \ten_choice_one_0_datasix_[1] , \ten_choice_one_0_datasix_[0] })
        , .dataseven({\ten_choice_one_0_dataseven_[11] , 
        \ten_choice_one_0_dataseven_[10] , 
        \ten_choice_one_0_dataseven_[9] , 
        \ten_choice_one_0_dataseven_[8] , 
        \ten_choice_one_0_dataseven_[7] , 
        \ten_choice_one_0_dataseven_[6] , 
        \ten_choice_one_0_dataseven_[5] , 
        \ten_choice_one_0_dataseven_[4] , 
        \ten_choice_one_0_dataseven_[3] , 
        \ten_choice_one_0_dataseven_[2] , 
        \ten_choice_one_0_dataseven_[1] , 
        \ten_choice_one_0_dataseven_[0] }), .dataeight({
        \ten_choice_one_0_dataeight_[11] , 
        \ten_choice_one_0_dataeight_[10] , 
        \ten_choice_one_0_dataeight_[9] , 
        \ten_choice_one_0_dataeight_[8] , 
        \ten_choice_one_0_dataeight_[7] , 
        \ten_choice_one_0_dataeight_[6] , 
        \ten_choice_one_0_dataeight_[5] , 
        \ten_choice_one_0_dataeight_[4] , 
        \ten_choice_one_0_dataeight_[3] , 
        \ten_choice_one_0_dataeight_[2] , 
        \ten_choice_one_0_dataeight_[1] , 
        \ten_choice_one_0_dataeight_[0] }), .datain({s_ADC[11], 
        s_ADC[10], s_ADC[9], s_ADC[8], s_ADC[7], s_ADC[6], s_ADC[5], 
        s_ADC[4], s_ADC[3], s_ADC[2], s_ADC[1], s_ADC[0]}));
    
endmodule
