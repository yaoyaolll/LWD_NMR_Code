library verilog;
use verilog.vl_types.all;
entity DUMP_OFF_DUMP_OFF_0 is
    port(
        bri_dump_sw_0_dumpoff_ctr: in     vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic;
        DUMP_OFF_0_dump_off: out    vl_logic;
        GLA             : in     vl_logic
    );
end DUMP_OFF_DUMP_OFF_0;
