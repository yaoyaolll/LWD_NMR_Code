library verilog;
use verilog.vl_types.all;
entity off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_4 is
    port(
        count_7         : out    vl_logic_vector(4 downto 0);
        GLA             : in     vl_logic;
        state1ms_choice_0_reset_out: in     vl_logic;
        off_on_state_1_state_over: in     vl_logic;
        dump_state_0_on_start: in     vl_logic
    );
end off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_4;
