library verilog;
use verilog.vl_types.all;
entity rst_n_module is
    port(
        rst_n_module_VCC: in     vl_logic;
        INV_0_Y         : in     vl_logic;
        GLA             : in     vl_logic;
        net_27          : out    vl_logic
    );
end rst_n_module;
