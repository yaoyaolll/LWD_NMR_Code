library verilog;
use verilog.vl_types.all;
entity off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1 is
    port(
        i_3             : in     vl_logic_vector(1 downto 0);
        GLA             : in     vl_logic;
        DUMP_OFF_0_dump_off: out    vl_logic;
        off_on_state_0_state_over: out    vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic
    );
end off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1;
