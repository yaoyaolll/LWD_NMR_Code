library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_3 is
    port(
        addresult_RNIDU3E: out    vl_logic_vector(4 downto 4);
        signal_data_iv_0_0_6: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_6_0: out    vl_logic;
        signal_data_iv_0_6_3: out    vl_logic;
        signal_data_iv_0_6_2: out    vl_logic;
        un1_n_s_change_0_1: in     vl_logic_vector(3 downto 0);
        un1_ten_choice_one_0_1_0: in     vl_logic;
        un1_ten_choice_one_0_1_2: in     vl_logic;
        un1_ten_choice_one_0_1_10: in     vl_logic;
        un1_ten_choice_one_0_1_5: in     vl_logic;
        un1_ten_choice_one_0_1_9: in     vl_logic;
        un1_ten_choice_one_0_1_7: in     vl_logic;
        un1_ten_choice_one_0_1_1: in     vl_logic;
        un1_ten_choice_one_0_1_8: in     vl_logic;
        un1_ten_choice_one_0_1_4: in     vl_logic;
        un1_ten_choice_one_0_1_6: in     vl_logic;
        un1_ten_choice_one_0_1_11: in     vl_logic;
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_249           : in     vl_logic;
        N_224           : out    vl_logic;
        N_91            : out    vl_logic;
        N_107           : out    vl_logic;
        N_192           : out    vl_logic;
        N_208           : out    vl_logic;
        N_251           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_241           : out    vl_logic;
        N_179           : out    vl_logic;
        N_171           : out    vl_logic;
        N_155           : out    vl_logic;
        N_147           : out    vl_logic;
        N_139           : out    vl_logic;
        N_131           : out    vl_logic;
        N_123           : out    vl_logic;
        N_115           : out    vl_logic;
        N_254           : in     vl_logic;
        N_99            : out    vl_logic;
        N_194           : in     vl_logic;
        N_243           : in     vl_logic;
        N_210_0         : in     vl_logic;
        N_226           : in     vl_logic;
        N_273           : in     vl_logic;
        N_213           : in     vl_logic;
        N_210           : in     vl_logic;
        N_216           : in     vl_logic
    );
end add_reg_add_reg_2_3;
