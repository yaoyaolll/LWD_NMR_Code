library verilog;
use verilog.vl_types.all;
entity off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_1 is
    port(
        count_6         : out    vl_logic_vector(4 downto 0);
        GLA             : in     vl_logic;
        OR2_2_Y         : in     vl_logic;
        off_on_state_0_state_over: in     vl_logic;
        OR2_1_Y         : in     vl_logic
    );
end off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_1;
