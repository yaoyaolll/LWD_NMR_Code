library verilog;
use verilog.vl_types.all;
entity qq_state_qq_state_0 is
    port(
        i_1             : in     vl_logic_vector(3 downto 1);
        i_2             : in     vl_logic_vector(0 downto 0);
        GLA             : in     vl_logic;
        Q1Q8_c          : out    vl_logic;
        qq_state_0_stateover: out    vl_logic;
        Q3Q6_c          : out    vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic
    );
end qq_state_qq_state_0;
