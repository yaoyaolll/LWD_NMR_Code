library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_1 is
    port(
        addresult_RNI8MQ7: out    vl_logic_vector(14 downto 14);
        addresult_RNIFE5C: in     vl_logic_vector(10 downto 10);
        signal_data_0_iv_i_2: in     vl_logic_vector(11 downto 4);
        addresult_RNIBOIB: in     vl_logic_vector(5 downto 5);
        signal_data_0_iv_i_5: out    vl_logic_vector(11 downto 4);
        signal_data_iv_0_0_3: in     vl_logic_vector(1 downto 1);
        signal_data_iv_0_0_9: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_3_0: in     vl_logic;
        signal_data_iv_0_3_3: in     vl_logic;
        signal_data_iv_0_3_2: in     vl_logic;
        signal_data_iv_0_9_0: out    vl_logic;
        signal_data_iv_0_9_3: out    vl_logic;
        signal_data_iv_0_9_2: out    vl_logic;
        un1_n_s_change_0_1: in     vl_logic_vector(4 downto 0);
        un1_ten_choice_one_0_5: in     vl_logic_vector(11 downto 0);
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_216           : out    vl_logic;
        N_249           : in     vl_logic;
        N_184           : out    vl_logic;
        N_200           : out    vl_logic;
        N_255           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_233           : out    vl_logic;
        N_262           : in     vl_logic;
        N_111           : out    vl_logic;
        N_95            : out    vl_logic;
        N_250           : in     vl_logic;
        N_87            : out    vl_logic;
        N_210           : in     vl_logic;
        N_214           : in     vl_logic;
        N_186           : in     vl_logic;
        N_174           : in     vl_logic;
        N_158           : in     vl_logic;
        N_134           : in     vl_logic;
        N_126           : in     vl_logic;
        N_118           : in     vl_logic;
        N_150           : in     vl_logic;
        N_235           : in     vl_logic;
        N_202           : in     vl_logic;
        N_218           : in     vl_logic;
        N_223           : in     vl_logic
    );
end add_reg_add_reg_2_1;
