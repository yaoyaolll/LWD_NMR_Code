library verilog;
use verilog.vl_types.all;
entity off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_2 is
    port(
        un1_off_on_timer_0: out    vl_logic_vector(4 downto 0);
        GLA             : in     vl_logic;
        nsctrl_choice_0_dumponoff_rst: in     vl_logic;
        off_on_state_0_state_over: in     vl_logic;
        nsctrl_choice_0_dumpoff_ctr: in     vl_logic
    );
end off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_2;
