library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_5 is
    port(
        s_addchoice     : in     vl_logic_vector(0 downto 0);
        signal_data_iv_0_0_13: in     vl_logic_vector(1 downto 1);
        signal_data_en  : in     vl_logic_vector(9 downto 9);
        signal_data_iv_0_13_2: in     vl_logic;
        signal_data_iv_0_13_3: in     vl_logic;
        signal_data_iv_0_13_0: in     vl_logic;
        un1_signal_acq_0: out    vl_logic_vector(3 downto 0);
        dataeight_0_a2_0_0: in     vl_logic_vector(0 downto 0);
        signal_data_0_iv_i_0: out    vl_logic_vector(11 downto 4);
        signal_data_iv_0_0_9: in     vl_logic_vector(1 downto 1);
        signal_data_iv_0_0_1: in     vl_logic_vector(1 downto 1);
        signal_data_iv_0_9_0: in     vl_logic;
        signal_data_iv_0_9_3: in     vl_logic;
        signal_data_iv_0_9_2: in     vl_logic;
        signal_data_iv_0_1_0: in     vl_logic;
        signal_data_iv_0_1_3: in     vl_logic;
        signal_data_iv_0_1_2: in     vl_logic;
        addresult_14    : out    vl_logic;
        addresult_13    : out    vl_logic;
        addresult_15    : out    vl_logic;
        addresult_12    : out    vl_logic;
        un1_ten_choice_one_0_7_2: in     vl_logic;
        un1_ten_choice_one_0_7_3: in     vl_logic;
        un1_ten_choice_one_0_7_5: in     vl_logic;
        un1_ten_choice_one_0_7_6: in     vl_logic;
        un1_ten_choice_one_0_7_7: in     vl_logic;
        un1_ten_choice_one_0_7_8: in     vl_logic;
        un1_ten_choice_one_0_7_9: in     vl_logic;
        un1_ten_choice_one_0_7_10: in     vl_logic;
        un1_ten_choice_one_0_7_11: in     vl_logic;
        un1_ten_choice_one_0_7_0: in     vl_logic;
        un1_n_s_change_0_1: in     vl_logic_vector(4 downto 0);
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_228           : out    vl_logic;
        N_245           : out    vl_logic;
        N_196           : out    vl_logic;
        G_1_0_a2_0      : in     vl_logic;
        N_212           : out    vl_logic;
        N_213           : in     vl_logic;
        N_182           : in     vl_logic;
        N_33            : in     vl_logic;
        N_256           : in     vl_logic;
        N_231           : in     vl_logic;
        N_198           : in     vl_logic;
        N_214           : in     vl_logic;
        N_267           : in     vl_logic;
        N_220           : in     vl_logic
    );
end add_reg_add_reg_2_5;
