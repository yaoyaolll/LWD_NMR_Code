library verilog;
use verilog.vl_types.all;
entity DUMP_OFF_DUMP_OFF_0_1 is
    port(
        nsctrl_choice_0_dumpoff_ctr: in     vl_logic;
        nsctrl_choice_0_dumponoff_rst: in     vl_logic;
        DUMP_OFF_1_dump_off: out    vl_logic;
        GLA             : in     vl_logic
    );
end DUMP_OFF_DUMP_OFF_0_1;
