library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_4 is
    port(
        un1_n_s_change_0_1: in     vl_logic_vector(2 downto 0);
        signal_data_0_iv_i_5: in     vl_logic_vector(11 downto 4);
        signal_data_0_iv_i_3: in     vl_logic_vector(11 downto 4);
        signal_data_0_iv_i_0: in     vl_logic_vector(11 downto 4);
        signal_data_iv_0_0_10: in     vl_logic_vector(1 downto 1);
        signal_data_iv_0_0_6: in     vl_logic_vector(1 downto 1);
        signal_data_iv_0_0_13: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_10_0: in     vl_logic;
        signal_data_iv_0_10_3: in     vl_logic;
        signal_data_iv_0_10_2: in     vl_logic;
        signal_data_iv_0_6_0: in     vl_logic;
        signal_data_iv_0_6_3: in     vl_logic;
        signal_data_iv_0_6_2: in     vl_logic;
        signal_data_iv_0_13_0: out    vl_logic;
        signal_data_iv_0_13_3: out    vl_logic;
        signal_data_iv_0_13_2: out    vl_logic;
        un1_ten_choice_one_0: in     vl_logic_vector(11 downto 0);
        addresult_4_10  : out    vl_logic;
        addresult_4_8   : out    vl_logic;
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_226           : out    vl_logic;
        N_249           : in     vl_logic;
        N_194           : out    vl_logic;
        N_210           : out    vl_logic;
        N_254           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_243           : out    vl_logic;
        N_108           : out    vl_logic;
        N_92            : out    vl_logic;
        N_222           : in     vl_logic;
        N_25_i_0        : out    vl_logic;
        N_20_i_0        : out    vl_logic;
        N_12_i_0        : out    vl_logic;
        N_14_i_0        : out    vl_logic;
        N_16_i_0        : out    vl_logic;
        N_18_i_0        : out    vl_logic;
        N_22_i_0        : out    vl_logic;
        N_27_i_0        : out    vl_logic;
        N_196           : in     vl_logic;
        N_39            : in     vl_logic;
        N_245           : in     vl_logic;
        N_212           : in     vl_logic;
        N_228           : in     vl_logic;
        N_271           : in     vl_logic
    );
end add_reg_add_reg_2_4;
