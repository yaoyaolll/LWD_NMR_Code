library verilog;
use verilog.vl_types.all;
entity qq_timer_qq_timer_0 is
    port(
        count_1         : out    vl_logic_vector(4 downto 0);
        GLA             : in     vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic;
        up              : in     vl_logic;
        qq_state_0_stateover: in     vl_logic
    );
end qq_timer_qq_timer_0;
