library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_6 is
    port(
        addresult_RNIJE5C: out    vl_logic_vector(14 downto 14);
        addresult_RNIFE5C: out    vl_logic_vector(10 downto 10);
        addresult_RNIBOIB: out    vl_logic_vector(5 downto 5);
        addresult_0_15  : out    vl_logic;
        addresult_0_13  : out    vl_logic;
        signal_data_iv_0_0_1: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_1_0: out    vl_logic;
        signal_data_iv_0_1_3: out    vl_logic;
        signal_data_iv_0_1_2: out    vl_logic;
        un1_n_s_change_0_1: in     vl_logic_vector(2 downto 0);
        un1_ten_choice_one_0_6: in     vl_logic_vector(11 downto 1);
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_214           : out    vl_logic;
        N_182           : out    vl_logic;
        N_221           : in     vl_logic;
        N_249           : in     vl_logic;
        N_198           : out    vl_logic;
        N_256           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_231           : out    vl_logic;
        N_174           : out    vl_logic;
        N_158           : out    vl_logic;
        N_150           : out    vl_logic;
        N_134           : out    vl_logic;
        N_126           : out    vl_logic;
        N_118           : out    vl_logic;
        N_255           : in     vl_logic;
        N_86            : out    vl_logic;
        N_210           : in     vl_logic;
        N_212           : in     vl_logic;
        N_184           : in     vl_logic;
        N_233           : in     vl_logic;
        N_200           : in     vl_logic;
        N_216           : in     vl_logic;
        N_270           : in     vl_logic
    );
end add_reg_add_reg_2_6;
