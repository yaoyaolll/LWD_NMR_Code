library verilog;
use verilog.vl_types.all;
entity add_reg_6 is
    port(
        dataone_0_a2_9  : in     vl_logic;
        dataone_0_a2_0  : in     vl_logic;
        ADC_c_3         : in     vl_logic;
        ADC_c_0_d0      : in     vl_logic;
        ADC_c_9         : in     vl_logic;
        ADC_c_5         : in     vl_logic;
        ADC_c_6         : in     vl_logic;
        ADC_c_8         : in     vl_logic;
        ADC_c_7         : in     vl_logic;
        ADC_c_4         : in     vl_logic;
        ADC_c_0_5       : in     vl_logic;
        ADC_c_0_0       : in     vl_logic;
        ADC_c_0_3       : in     vl_logic;
        ADC_c_0_4       : in     vl_logic;
        ADC_c_0_2       : in     vl_logic;
        ADC_c_0_6       : in     vl_logic;
        un1_ten_choice_one_0_0: in     vl_logic;
        un1_ten_choice_one_0_6: in     vl_logic;
        un1_ten_choice_one_0_9: in     vl_logic;
        addresult_7     : out    vl_logic_vector(31 downto 0);
        reset_c         : in     vl_logic;
        AND2_2_Y        : in     vl_logic;
        N_274           : in     vl_logic;
        ADD_32x32_fast_I169_Y_0_o2_5_m12_i_a7_3_0: in     vl_logic;
        N_264           : in     vl_logic;
        ADD_32x32_fast_I169_Y_0_o2_5_N_21: in     vl_logic;
        N_261           : in     vl_logic;
        N_274_0         : in     vl_logic
    );
end add_reg_6;
