library verilog;
use verilog.vl_types.all;
entity ten_choice_one is
    port(
        un1_ten_choice_one_0_7_0: out    vl_logic;
        un1_ten_choice_one_0_7_2: out    vl_logic;
        un1_ten_choice_one_0_7_11: out    vl_logic;
        un1_ten_choice_one_0_7_10: out    vl_logic;
        un1_ten_choice_one_0_7_9: out    vl_logic;
        un1_ten_choice_one_0_7_8: out    vl_logic;
        un1_ten_choice_one_0_7_7: out    vl_logic;
        un1_ten_choice_one_0_7_6: out    vl_logic;
        un1_ten_choice_one_0_7_5: out    vl_logic;
        un1_ten_choice_one_0_7_3: out    vl_logic;
        un1_ten_choice_one_0_4_3: out    vl_logic;
        un1_ten_choice_one_0_4_1: out    vl_logic;
        un1_ten_choice_one_0_4_0: out    vl_logic;
        un1_ten_choice_one_0_4_11: out    vl_logic;
        un1_ten_choice_one_0_4_10: out    vl_logic;
        un1_ten_choice_one_0_4_9: out    vl_logic;
        un1_ten_choice_one_0_4_8: out    vl_logic;
        un1_ten_choice_one_0_4_7: out    vl_logic;
        un1_ten_choice_one_0_4_6: out    vl_logic;
        un1_ten_choice_one_0_4_5: out    vl_logic;
        un1_ten_choice_one_0_4_4: out    vl_logic;
        un1_ten_choice_one_0_3_1: out    vl_logic;
        un1_ten_choice_one_0_3_0: out    vl_logic;
        un1_ten_choice_one_0_3_10: out    vl_logic;
        un1_ten_choice_one_0_3_11: out    vl_logic;
        un1_ten_choice_one_0_3_9: out    vl_logic;
        un1_ten_choice_one_0_3_8: out    vl_logic;
        un1_ten_choice_one_0_3_7: out    vl_logic;
        un1_ten_choice_one_0_3_6: out    vl_logic;
        un1_ten_choice_one_0_3_5: out    vl_logic;
        un1_ten_choice_one_0_3_4: out    vl_logic;
        un1_ten_choice_one_0_3_3: out    vl_logic;
        un1_ten_choice_one_0: out    vl_logic_vector(11 downto 0);
        un1_ten_choice_one_0_6: out    vl_logic_vector(11 downto 1);
        un1_ten_choice_one_0_5: out    vl_logic_vector(11 downto 0);
        un1_ten_choice_one_0_1_2: out    vl_logic;
        un1_ten_choice_one_0_1_1: out    vl_logic;
        un1_ten_choice_one_0_1_0: out    vl_logic;
        un1_ten_choice_one_0_1_8: out    vl_logic;
        un1_ten_choice_one_0_1_10: out    vl_logic;
        un1_ten_choice_one_0_1_11: out    vl_logic;
        un1_ten_choice_one_0_1_9: out    vl_logic;
        un1_ten_choice_one_0_1_7: out    vl_logic;
        un1_ten_choice_one_0_1_6: out    vl_logic;
        un1_ten_choice_one_0_1_5: out    vl_logic;
        un1_ten_choice_one_0_1_4: out    vl_logic;
        addrout         : in     vl_logic_vector(3 downto 0);
        dataeight_0_a2_0_0: out    vl_logic_vector(0 downto 0);
        un1_n_s_change_0_1: in     vl_logic_vector(11 downto 0);
        un1_ten_choice_one_0_2_0: out    vl_logic;
        un1_ten_choice_one_0_2_10: out    vl_logic;
        un1_ten_choice_one_0_2_9: out    vl_logic;
        un1_ten_choice_one_0_2_8: out    vl_logic;
        un1_ten_choice_one_0_2_7: out    vl_logic;
        un1_ten_choice_one_0_2_6: out    vl_logic;
        un1_ten_choice_one_0_2_5: out    vl_logic;
        un1_ten_choice_one_0_2_4: out    vl_logic;
        un1_ten_choice_one_0_2_3: out    vl_logic;
        un1_ten_choice_one_0_2_2: out    vl_logic;
        N_214           : out    vl_logic;
        N_212           : out    vl_logic;
        N_211           : out    vl_logic;
        N_217           : out    vl_logic;
        N_219           : out    vl_logic;
        N_222           : out    vl_logic;
        N_221           : out    vl_logic;
        N_223           : out    vl_logic;
        N_224           : out    vl_logic;
        N_216           : out    vl_logic;
        N_213           : out    vl_logic;
        N_220           : out    vl_logic;
        N_210           : out    vl_logic;
        N_215           : out    vl_logic
    );
end ten_choice_one;
