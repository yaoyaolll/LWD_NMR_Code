library verilog;
use verilog.vl_types.all;
entity qq_state_qq_state_0_1 is
    port(
        i               : in     vl_logic_vector(3 downto 1);
        i_0             : in     vl_logic_vector(0 downto 0);
        GLA             : in     vl_logic;
        Q2Q7_c          : out    vl_logic;
        qq_state_1_stateover: out    vl_logic;
        Q4Q5_c          : out    vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic
    );
end qq_state_qq_state_0_1;
