library verilog;
use verilog.vl_types.all;
entity off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_1 is
    port(
        i_5             : in     vl_logic_vector(1 downto 1);
        i_6             : in     vl_logic_vector(0 downto 0);
        GLA             : in     vl_logic;
        off_on_state_0_state_over: out    vl_logic;
        DUMP_ON_0_dump_on: out    vl_logic;
        OR2_2_Y         : in     vl_logic
    );
end off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_1;
