library verilog;
use verilog.vl_types.all;
entity NMR_TOP is
    port(
        zcs2            : in     vl_logic;
        xwe             : in     vl_logic;
        ddsfqud         : out    vl_logic;
        ddsreset        : out    vl_logic;
        ddswclk         : out    vl_logic;
        cal_out         : out    vl_logic;
        ddsdata         : out    vl_logic;
        OCX40MHz        : in     vl_logic;
        ddsclkout       : in     vl_logic;
        interupt        : out    vl_logic;
        rt_sw           : out    vl_logic;
        soft_dump       : out    vl_logic;
        sw_acq1         : out    vl_logic;
        sw_acq2         : out    vl_logic;
        dumpon          : out    vl_logic;
        dumpoff         : out    vl_logic;
        Q1Q8            : out    vl_logic;
        Q3Q6            : out    vl_logic;
        Q4Q5            : out    vl_logic;
        Q2Q7            : out    vl_logic;
        calcuinter      : out    vl_logic;
        tri_ctrl        : in     vl_logic;
        sigtimeup       : out    vl_logic;
        k1              : out    vl_logic;
        k2              : out    vl_logic;
        gpio            : in     vl_logic;
        pulse_start     : out    vl_logic;
        pd_pulse_en     : out    vl_logic;
        XRD             : in     vl_logic;
        Acq_clk         : out    vl_logic;
        sd_acq_en       : out    vl_logic;
        s_acq180        : out    vl_logic;
        GLA             : out    vl_logic;
        xa              : in     vl_logic_vector(18 downto 0);
        xd              : inout  vl_logic_vector(15 downto 0);
        relayclose_on   : out    vl_logic_vector(15 downto 0);
        ADC             : in     vl_logic_vector(11 downto 0)
    );
end NMR_TOP;
