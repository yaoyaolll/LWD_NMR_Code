library verilog;
use verilog.vl_types.all;
entity off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_2 is
    port(
        un1_off_on_coder_0: in     vl_logic_vector(1 downto 0);
        GLA             : in     vl_logic;
        DUMP_OFF_1_dump_off: out    vl_logic;
        off_on_state_0_state_over: out    vl_logic;
        nsctrl_choice_0_dumponoff_rst: in     vl_logic
    );
end off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_2;
