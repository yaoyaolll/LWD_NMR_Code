library verilog;
use verilog.vl_types.all;
entity dump_sustain_timer_tb is
end dump_sustain_timer_tb;
