library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_2 is
    port(
        addresult_RNIVJME: out    vl_logic_vector(4 downto 4);
        un1_n_s_change_0_1: in     vl_logic_vector(2 downto 0);
        un1_ten_choice_one_0_3_0: in     vl_logic;
        un1_ten_choice_one_0_3_1: in     vl_logic;
        un1_ten_choice_one_0_3_3: in     vl_logic;
        un1_ten_choice_one_0_3_10: in     vl_logic;
        un1_ten_choice_one_0_3_4: in     vl_logic;
        un1_ten_choice_one_0_3_6: in     vl_logic;
        un1_ten_choice_one_0_3_7: in     vl_logic;
        un1_ten_choice_one_0_3_8: in     vl_logic;
        un1_ten_choice_one_0_3_9: in     vl_logic;
        un1_ten_choice_one_0_3_11: in     vl_logic;
        un1_ten_choice_one_0_3_5: in     vl_logic;
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_249           : in     vl_logic;
        N_220           : out    vl_logic;
        N_221           : out    vl_logic;
        N_205           : out    vl_logic;
        N_89            : out    vl_logic;
        N_105           : out    vl_logic;
        N_204           : out    vl_logic;
        N_189           : out    vl_logic;
        N_266           : in     vl_logic;
        N_238           : out    vl_logic;
        N_237           : out    vl_logic;
        N_253           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_188           : out    vl_logic;
        N_177           : out    vl_logic;
        N_169           : out    vl_logic;
        N_153           : out    vl_logic;
        N_145           : out    vl_logic;
        N_137           : out    vl_logic;
        N_129           : out    vl_logic;
        N_121           : out    vl_logic;
        N_113           : out    vl_logic;
        N_252           : in     vl_logic;
        N_97            : out    vl_logic;
        N_219           : in     vl_logic
    );
end add_reg_add_reg_2_2;
