`timescale 1 ns/100 ps
// Version: 9.1 9.1.0.18


module state1ms_choice(
       state1ms_choice_0_bri_cycle,
       state1ms_choice_0_dump_start,
       bri_div_start_0,
       state1ms_choice_0_reset_out,
       rt_sw_c,
       GLA,
       soft_dump_c,
       state_1ms_0_soft_dump,
       soft_dump_net_1,
       state_1ms_0_rt_sw,
       rt_sw_net_1,
       state_1ms_0_reset_out,
       bri_dump_sw_0_reset_out_0,
       state_1ms_0_pluse_start,
       bri_dump_sw_0_off_test,
       state_1ms_0_dump_start,
       bri_dump_sw_0_dump_start,
       top_code_0_state_1ms_start,
       state_1ms_0_bri_cycle,
       PLUSE_0_bri_cycle,
       net_27
    );
output state1ms_choice_0_bri_cycle;
output state1ms_choice_0_dump_start;
output bri_div_start_0;
output state1ms_choice_0_reset_out;
output rt_sw_c;
input  GLA;
output soft_dump_c;
input  state_1ms_0_soft_dump;
input  soft_dump_net_1;
input  state_1ms_0_rt_sw;
input  rt_sw_net_1;
input  state_1ms_0_reset_out;
input  bri_dump_sw_0_reset_out_0;
input  state_1ms_0_pluse_start;
input  bri_dump_sw_0_off_test;
input  state_1ms_0_dump_start;
input  bri_dump_sw_0_dump_start;
input  top_code_0_state_1ms_start;
input  state_1ms_0_bri_cycle;
input  PLUSE_0_bri_cycle;
input  net_27;

    wire reset_out_RNO_net_1, reset_out_5, pluse_start_RNO_net_1, 
        pluse_start_5, dump_start_RNO_net_1, dump_start_5, 
        bri_cycle_RNO_net_1, bri_cycle_5, rt_sw_4, soft_dump_4, GND, 
        VCC, GND_0, VCC_0;
    
    DFN1E1 rt_sw (.D(rt_sw_4), .CLK(GLA), .E(net_27), .Q(rt_sw_c));
    NOR2A reset_out_RNO (.A(net_27), .B(reset_out_5), .Y(
        reset_out_RNO_net_1));
    DFN1 dump_start (.D(dump_start_RNO_net_1), .CLK(GLA), .Q(
        state1ms_choice_0_dump_start));
    MX2 soft_dump_RNO (.A(soft_dump_net_1), .B(state_1ms_0_soft_dump), 
        .S(top_code_0_state_1ms_start), .Y(soft_dump_4));
    GND GND_i_0 (.Y(GND_0));
    MX2C pluse_start_RNO_0 (.A(bri_dump_sw_0_off_test), .B(
        state_1ms_0_pluse_start), .S(top_code_0_state_1ms_start), .Y(
        pluse_start_5));
    VCC VCC_i (.Y(VCC));
    NOR2A bri_cycle_RNO (.A(net_27), .B(bri_cycle_5), .Y(
        bri_cycle_RNO_net_1));
    GND GND_i (.Y(GND));
    MX2C dump_start_RNO_0 (.A(bri_dump_sw_0_dump_start), .B(
        state_1ms_0_dump_start), .S(top_code_0_state_1ms_start), .Y(
        dump_start_5));
    MX2C bri_cycle_RNO_0 (.A(PLUSE_0_bri_cycle), .B(
        state_1ms_0_bri_cycle), .S(top_code_0_state_1ms_start), .Y(
        bri_cycle_5));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1E1 soft_dump (.D(soft_dump_4), .CLK(GLA), .E(net_27), .Q(
        soft_dump_c));
    MX2 rt_sw_RNO (.A(rt_sw_net_1), .B(state_1ms_0_rt_sw), .S(
        top_code_0_state_1ms_start), .Y(rt_sw_4));
    MX2C reset_out_RNO_0 (.A(bri_dump_sw_0_reset_out_0), .B(
        state_1ms_0_reset_out), .S(top_code_0_state_1ms_start), .Y(
        reset_out_5));
    DFN1 pluse_start (.D(pluse_start_RNO_net_1), .CLK(GLA), .Q(
        bri_div_start_0));
    NOR2A dump_start_RNO (.A(net_27), .B(dump_start_5), .Y(
        dump_start_RNO_net_1));
    NOR2A pluse_start_RNO (.A(net_27), .B(pluse_start_5), .Y(
        pluse_start_RNO_net_1));
    DFN1 reset_out (.D(reset_out_RNO_net_1), .CLK(GLA), .Q(
        state1ms_choice_0_reset_out));
    DFN1 bri_cycle (.D(bri_cycle_RNO_net_1), .CLK(GLA), .Q(
        state1ms_choice_0_bri_cycle));
    
endmodule


module top_code(
       plusedata,
       s_acqnum_0,
       s_addchoice,
       s_periodnum,
       scalechoice,
       scaledatain,
       scaleddsdiv,
       scandata,
       sd_sacq_choice,
       sd_sacq_data,
       sigtimedata,
       state_1ms_data,
       state_1ms_lc,
       bri_datain,
       cal_data,
       change,
       dds_configdata,
       dump_cho,
       dumpdata,
       halfdata,
       n_acqnum,
       n_divnum,
       noisedata,
       pd_pluse_choice,
       pd_pluse_data,
       un1_GPMI_0_1,
       relayclose_on_c,
       xa_c_0_0,
       xa_c_0_7,
       xa_c,
       un1_GPMI_0_1_0,
       un1_top_code_0_3_0,
       net_33,
       top_code_0_noise_rst,
       top_code_0_bridge_load,
       top_code_0_scale_start,
       top_code_0_pn_change,
       top_code_0_scanload,
       top_code_0_acqclken,
       top_code_0_state_1ms_rst_n,
       top_code_0_scaleload,
       top_code_0_scan_start,
       top_code_0_n_load,
       top_code_0_n_rd_en,
       top_code_0_n_s_ctrl,
       top_code_0_RAM_Rd_rst,
       top_code_0_noise_start,
       top_code_0_dds_choice,
       top_code_0_dumpload,
       top_code_0_pluseload,
       top_code_0_scanchoice,
       top_code_0_pluse_scale,
       top_code_0_state_1ms_load,
       top_code_0_sd_sacq_load,
       top_code_0_pd_pluse_load,
       top_code_0_nstateload,
       top_code_0_pluse_lc,
       top_code_0_sigrst,
       top_code_0_s_load,
       top_code_0_cal_load,
       top_code_0_nstatechoice,
       top_code_0_pluse_noise_ctrl,
       top_code_0_dump_sustain,
       k1_c,
       k2_c,
       top_code_0_pluse_rst,
       top_code_0_pluse_str,
       top_code_0_state_1ms_start,
       GPMI_0_code_en,
       top_code_0_scale_rst,
       top_code_0_dds_load,
       top_code_0_n_s_ctrl_0,
       top_code_0_n_s_ctrl_1,
       top_code_0_state_1ms_rst_n_0,
       net_27,
       top_code_0_bridge_load_0,
       net_33_0,
       top_code_0_pluse_rst_0,
       GLA,
       top_code_0_noise_rst_0
    );
output [15:0] plusedata;
output [15:0] s_acqnum_0;
output [4:0] s_addchoice;
output [3:0] s_periodnum;
output [4:0] scalechoice;
output [15:0] scaledatain;
output [5:0] scaleddsdiv;
output [15:0] scandata;
output [3:0] sd_sacq_choice;
output [15:0] sd_sacq_data;
output [15:0] sigtimedata;
output [15:0] state_1ms_data;
output [3:0] state_1ms_lc;
output [15:0] bri_datain;
output [5:0] cal_data;
output [1:0] change;
output [15:0] dds_configdata;
output [2:0] dump_cho;
output [11:0] dumpdata;
output [7:0] halfdata;
output [11:0] n_acqnum;
output [9:0] n_divnum;
output [15:0] noisedata;
output [3:0] pd_pluse_choice;
output [15:0] pd_pluse_data;
input  [15:0] un1_GPMI_0_1;
output [15:0] relayclose_on_c;
input  xa_c_0_0;
input  xa_c_0_7;
input  [18:0] xa_c;
input  [2:0] un1_GPMI_0_1_0;
output [1:0] un1_top_code_0_3_0;
output net_33;
output top_code_0_noise_rst;
output top_code_0_bridge_load;
output top_code_0_scale_start;
output top_code_0_pn_change;
output top_code_0_scanload;
output top_code_0_acqclken;
output top_code_0_state_1ms_rst_n;
output top_code_0_scaleload;
output top_code_0_scan_start;
output top_code_0_n_load;
output top_code_0_n_rd_en;
output top_code_0_n_s_ctrl;
output top_code_0_RAM_Rd_rst;
output top_code_0_noise_start;
output top_code_0_dds_choice;
output top_code_0_dumpload;
output top_code_0_pluseload;
output top_code_0_scanchoice;
output top_code_0_pluse_scale;
output top_code_0_state_1ms_load;
output top_code_0_sd_sacq_load;
output top_code_0_pd_pluse_load;
output top_code_0_nstateload;
output top_code_0_pluse_lc;
output top_code_0_sigrst;
output top_code_0_s_load;
output top_code_0_cal_load;
output top_code_0_nstatechoice;
output top_code_0_pluse_noise_ctrl;
output top_code_0_dump_sustain;
output k1_c;
output k2_c;
output top_code_0_pluse_rst;
output top_code_0_pluse_str;
output top_code_0_state_1ms_start;
input  GPMI_0_code_en;
output top_code_0_scale_rst;
output top_code_0_dds_load;
output top_code_0_n_s_ctrl_0;
output top_code_0_n_s_ctrl_1;
output top_code_0_state_1ms_rst_n_0;
input  net_27;
output top_code_0_bridge_load_0;
output net_33_0;
output top_code_0_pluse_rst_0;
input  GLA;
output top_code_0_noise_rst_0;

    wire N_38, N_41, change_1_sqmuxa, N_43, N_181, N_225, n_s_ctrl_3, 
        dds_load_net_1, scale_rst_net_1, 
        state_1ms_data_1_sqmuxa_0_a2_0_net_1, 
        noisedata_1_sqmuxa_0_a2_1_net_1, N_280, N_122, 
        un1_state_1ms_rst_n113_45_i_a2_0_0, 
        scalechoice_1_sqmuxa_0_a2_0_a2_0_net_1, N_278, N_445, 
        un1_state_1ms_rst_n113_43_i_a2_2_0_net_1, N_232, 
        un1_state_1ms_rst_n113_44_i_a2_0_0, N_229, 
        scaleload_3_i_i_a2_0_0, scanload_3_i_a2_0_0, N_128, N_132, 
        pn_change_3_0_i_o2_0_net_1, pn_change_3_0_i_a2_0_0, 
        n_s_ctrl_3_0_a2_0_6_net_1, n_s_ctrl_3_0_a2_0_1_net_1, 
        n_s_ctrl_3_0_a2_0_0_net_1, n_s_ctrl_3_0_a2_0_5_net_1, 
        n_s_ctrl_3_0_a2_0_3_net_1, un1_xa_7_3, N_262, 
        scanchoice_3_i_a2_0_1, N_138, scanchoice_3_i_a2_0_0, 
        dds_choice_3_0_o2_1_net_1, cal_load_3_i_i_a2_0_0, N_277, 
        relayclose_on_1_sqmuxa_0_a2_2_a2_3_net_1, 
        relayclose_on_1_sqmuxa_0_a2_2_a2_2_net_1, N_297, 
        dds_choice_3_0_a2_0_2, N_125, dds_choice_3_0_a2_0_1, N_1559, 
        n_s_ctrl_3_0_o2_0, N_141, N_147, sigrst_3_i_a2_0_0, 
        un1_state_1ms_rst_n113_5_i_a2_0_a2_0, N_282, acqclken_3_0_o2_2, 
        N_121, acqclken_3_0_o2_1, N_260, N_272, 
        un1_state_1ms_rst_n113_28_i_a2_2_net_1, N_120_i, 
        un1_state_1ms_rst_n113_28_i_a2_1_net_1, N_136, 
        un1_state_1ms_rst_n113_35_i_a2_1, 
        un1_state_1ms_rst_n113_35_i_a2_0, N_233, 
        pluse_scale_3_0_a2_0_4, pluse_scale_3_0_a2_0_1, 
        pluse_scale_3_0_a2_0_0, pluse_scale_3_0_a2_0_2, N_158, N_264, 
        N_144_i_0, acqclken_3_0_a2_0_3, acqclken_3_0_a2_0_2, 
        N_220_1_i_0, N_150, pluse_scale_3_0_o2_1, N_134, 
        nstatechoice_3_0_i_o2_1_m1_e_2_net_1, 
        dumpload_3_i_i_o2_0_net_1, 
        nstatechoice_3_0_i_o2_1_m1_e_1_net_1, 
        acqclken_3_0_o2_0_0_1_net_1, acqclken_3_0_o2_0_0_0_net_1, 
        un1_state_1ms_rst_n113_41_i_a2_1_0, un1_xa_10_0_a2_0_a2_0, 
        un1_state_1ms_rst_n113_42_i_a2_1_0, un1_xa_131_3_1_net_1, 
        un1_xa_10, un1_xa_13, un1_xa_131_3_0_net_1, 
        un1_xa_131_2_0_a2_2_net_1, un1_xa_131_2_0_a2_1_net_1, un1_xa_4, 
        un1_xa_10_0_a2_0_a2_1_net_1, un1_xa_49_0_a2_1_net_1, N_315, 
        N_276, N_178, N_151, N_1554, N_191, N_352, N_190, un1_xa_49, 
        N_238, N_197, N_235, N_119, N_268, scandata_1_sqmuxa, N_288, 
        N_163_1, N_446, N_214, N_140, N_164, N_293, 
        s_addchoice_1_sqmuxa, N_299, N_228, N_458, plusedata_1_sqmuxa, 
        N_462, cal_data_1_sqmuxa, N_286, N_1395, n_acqnum_1_sqmuxa, 
        N_290, halfdata_1_sqmuxa, N_287, N_459, state_1ms_lc_1_sqmuxa, 
        N_451, s_periodnum_1_sqmuxa, sigtimedata_1_sqmuxa, 
        state_1ms_data_1_sqmuxa, N_341, dump_cho_1_sqmuxa, N_222, 
        N_411_1, N_156, N_1562, N_200, N_186_2, N_29, N_188, 
        noise_start_RNO_2_net_1, N_31_2, N_176, N_239, N_210, N_1558, 
        relayclose_on_1_sqmuxa, N_31, un1_state_1ms_rst_n113_42_i_0, 
        noisedata_1_sqmuxa, N_157, scalechoice_1_sqmuxa, N_209, 
        un1_xa_2, N_148, N_263, N_275, N_351_i, N_448, N_393, 
        un1_state_1ms_rst_n113_42_i_a2_1, 
        un1_state_1ms_rst_n113_43_i_a2_0_1, 
        un1_state_1ms_rst_n113_41_i_a2_1, 
        un1_state_1ms_rst_n113_43_i_a2_0, N_123, N_783, N_786, N_28, 
        N_790, N_791, N_163, N_792, N_793, N_1449, N_794, N_118, N_795, 
        N_796, N_803, N_804, N_806, N_807, N_808, N_809, N_810, N_355, 
        N_296, scaleddsdiv_1_sqmuxa, N_371, N_300, N_377, N_279, N_379, 
        N_294, N_395, N_292, N_396, N_295, N_408, N_309, 
        bri_datain_1_sqmuxa, pd_pluse_choice_1_sqmuxa, 
        sd_sacq_data_1_sqmuxa, n_divnum_1_sqmuxa, scaledatain_1_sqmuxa, 
        pd_pluse_data_1_sqmuxa, N_461, N_6, N_317, N_30, N_316, N_1542, 
        N_303, N_70, N_311, N_82, N_325, N_1543, N_106, N_1544, N_381, 
        N_179, N_319, N_201, N_310, N_203, N_327, N_192, N_160, N_215, 
        state_1ms_load_RNO_net_1, N_159, N_12, pluseload_3, N_1565, 
        pluse_scale_3, N_52, N_54, N_59, N_62, N_66, N_69, N_71, N_79, 
        N_81, N_83, N_87, N_93, N_95, dumpdata_1_sqmuxa, 
        sd_sacq_choice_1_sqmuxa_1, N_45, N_130, N_85, N_787, 
        dds_choice_3, N_124, N_269, N_789, un1_xa_30, N_223, N_101, 
        N_799, N_91, N_784, N_217, N_129, N_320, N_205, N_410, N_168, 
        N_386, dds_configdata_1_sqmuxa, s_acqnum_1_sqmuxa, 
        \relayclose_on_RNO[4]_net_1 , N_800, N_50, N_802, N_47, N_801, 
        N_175, N_390, N_99, N_798, N_97, N_797, N_73, N_811, N_56, 
        N_805, N_788, sd_sacq_choice_1_sqmuxa, N_89, N_785, acqclken_3, 
        N_219, N_1556_i_0, N_194_i, N_177, N_26, GND, VCC, GND_0, 
        VCC_0;
    
    DFN1E1 \dumpdata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[6]));
    DFN1E1 \s_periodnum[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        s_periodnum_1_sqmuxa), .Q(s_periodnum[0]));
    OA1B n_rd_en_RNO (.A(N_320), .B(top_code_0_n_rd_en), .C(N_386), .Y(
        N_168));
    DFN1E1 \sigtimedata[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[2]));
    MX2 \relayclose_on_RNO_0[0]  (.A(relayclose_on_c[0]), .B(
        un1_GPMI_0_1_0[0]), .S(relayclose_on_1_sqmuxa), .Y(N_796));
    DFN1E1 \dds_configdata[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[0]));
    DFN1E1 \scaledatain[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[3]));
    OR2 cal_load_3_i_i_o2_1 (.A(xa_c_0_7), .B(N_279), .Y(N_286));
    DFN1 \relayclose_on[9]  (.D(N_56), .CLK(GLA), .Q(
        relayclose_on_c[9]));
    DFN1E1 \plusedata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[3]));
    DFN1E1 \noisedata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[10]));
    MX2B state_1ms_start_RNO_0 (.A(top_code_0_state_1ms_start), .B(
        un1_xa_4), .S(N_1554), .Y(N_783));
    DFN1E1 \sd_sacq_data[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[0]));
    NOR3A pluse_lc_RNO_0 (.A(xa_c[7]), .B(N_277), .C(N_293), .Y(N_311));
    OR2 un1_xa_49_0_a2_1 (.A(xa_c_0_0), .B(xa_c[3]), .Y(
        un1_xa_49_0_a2_1_net_1));
    OR3 pluseload_RNO_1 (.A(N_1559), .B(N_238), .C(N_140), .Y(N_214));
    DFN1E1 \s_acqnum[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[12]));
    DFN1E1 \bri_datain[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[7]));
    DFN1E1 \pd_pluse_data[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[8]));
    DFN1E1 \s_periodnum[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        s_periodnum_1_sqmuxa), .Q(s_periodnum[3]));
    OR2A un1_xa_131_2_0_o2 (.A(xa_c[0]), .B(xa_c[2]), .Y(N_124));
    DFN1E1 \sigtimedata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[7]));
    OR2B un1_xa_131_2_0_o2_0 (.A(N_260), .B(N_121), .Y(N_122));
    OAI1 n_load_RNO_0 (.A(N_158), .B(N_290), .C(top_code_0_n_load), .Y(
        N_410));
    MX2 \relayclose_on_RNO_0[10]  (.A(relayclose_on_c[10]), .B(
        un1_GPMI_0_1[10]), .S(relayclose_on_1_sqmuxa), .Y(N_806));
    OR2 scan_start_RNO_4 (.A(un1_state_1ms_rst_n113_42_i_a2_1_0), .B(
        un1_xa_7_3), .Y(un1_state_1ms_rst_n113_42_i_a2_1));
    DFN1E1 \scandata[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[14]));
    MX2 scale_start_RNO_0 (.A(top_code_0_scale_start), .B(xa_c[0]), .S(
        N_26), .Y(N_785));
    OA1C pluse_noise_ctrl_RNO (.A(N_303), .B(N_300), .C(N_371), .Y(
        N_1542));
    DFN1E1 \plusedata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[7]));
    AO1A n_s_ctrl_RNIASSC5 (.A(N_235), .B(n_s_ctrl_3_0_a2_0_6_net_1), 
        .C(N_217), .Y(n_s_ctrl_3));
    DFN1E1 pluse_noise_ctrl (.D(N_1542), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pluse_noise_ctrl));
    MX2 \relayclose_on_RNO_0[13]  (.A(relayclose_on_c[13]), .B(
        un1_GPMI_0_1[13]), .S(relayclose_on_1_sqmuxa), .Y(N_809));
    DFN1E1 \scaledatain[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[0]));
    OR2A sd_sacq_choice_1_sqmuxa_0_a2_0_a2_1 (.A(N_287), .B(N_445), .Y(
        sd_sacq_choice_1_sqmuxa_1));
    CLKINT dds_load_RNIM024 (.A(dds_load_net_1), .Y(
        top_code_0_dds_load));
    OAI1 cal_load_RNO_1 (.A(N_280), .B(N_294), .C(top_code_0_cal_load), 
        .Y(N_379));
    DFN1E1 \halfdata[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[0]));
    OR2 scalechoice_1_sqmuxa_0_a2_0_a2_0 (.A(N_278), .B(N_445), .Y(
        scalechoice_1_sqmuxa_0_a2_0_a2_0_net_1));
    NOR2 s_acqnum_1_sqmuxa_0_a2_0_a2_0 (.A(N_446), .B(N_280), .Y(N_461)
        );
    DFN1E1 \dds_configdata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[7]));
    DFN1E1 \state_1ms_data[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[14]));
    NOR3 dumpdata_1_sqmuxa_0_a2_0_a2 (.A(N_276), .B(N_277), .C(
        sd_sacq_choice_1_sqmuxa_1), .Y(dumpdata_1_sqmuxa));
    DFN1E1 \s_acqnum[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[3]));
    DFN1E1 \cal_data[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[5]));
    OA1C scanchoice_RNO (.A(N_178), .B(top_code_0_scanchoice), .C(
        N_197), .Y(N_12));
    OR2A un1_xa_66_0_o2_0_i_o2 (.A(N_260), .B(xa_c[11]), .Y(N_262));
    MX2 pluse_rst_RNIM3QQ2 (.A(top_code_0_pluse_rst), .B(xa_c_0_0), .S(
        N_163), .Y(N_791));
    DFN1E1 \sd_sacq_data[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[4]));
    NOR2B pluse_str_RNO (.A(N_786), .B(net_27), .Y(N_87));
    DFN1E1 \pd_pluse_data[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[9]));
    DFN1E1 \scaledatain[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[6]));
    NOR2B \relayclose_on_RNO[15]  (.A(N_811), .B(net_27), .Y(N_73));
    DFN1E1 \sd_sacq_choice[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        sd_sacq_choice_1_sqmuxa), .Q(sd_sacq_choice[0]));
    NOR2B \relayclose_on_RNO[4]  (.A(N_800), .B(net_27), .Y(
        \relayclose_on_RNO[4]_net_1 ));
    NOR2B dump_sustain_RNO (.A(N_795), .B(net_27), .Y(N_79));
    DFN1E1 \bri_datain[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[12]));
    NOR3 cal_data_1_sqmuxa_0_a2_0_a2 (.A(N_286), .B(N_277), .C(N_445), 
        .Y(cal_data_1_sqmuxa));
    DFN1E1 \bri_datain[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[5]));
    OR2B un1_xa_10_0_a2_0_a2 (.A(un1_xa_10_0_a2_0_a2_1_net_1), .B(
        un1_xa_10_0_a2_0_a2_0), .Y(un1_xa_10));
    DFN1E1 \plusedata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[8]));
    DFN1E1 \n_divnum[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[7]));
    DFN1E1 \n_acqnum[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[6]));
    DFN1E1 \plusedata[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[0]));
    DFN1E1 \scandata[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[15]));
    OA1A scanload_RNO (.A(N_160), .B(scanload_3_i_a2_0_0), .C(N_194_i), 
        .Y(N_1556_i_0));
    NOR3B pd_pluse_load_RNO_0 (.A(N_292), .B(xa_c[7]), .C(N_272), .Y(
        N_319));
    DFN1E1 \plusedata[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[13]));
    NOR2B noise_start_RNO (.A(N_787), .B(net_27), .Y(N_85));
    NOR2 pluse_scale_RNO_4 (.A(xa_c[8]), .B(xa_c[9]), .Y(
        pluse_scale_3_0_a2_0_2));
    OA1B bridge_load_0_RNIJRSC5 (.A(N_276), .B(N_309), .C(N_396), .Y(
        N_181));
    DFN1E1 \s_addchoice[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        s_addchoice_1_sqmuxa), .Q(s_addchoice[4]));
    NOR2A sd_sacq_choice_1_sqmuxa_0_a2_0_o2 (.A(xa_c[4]), .B(xa_c[3]), 
        .Y(N_287));
    DFN1E1 \sigtimedata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[9]));
    NOR2B \relayclose_on_RNO[13]  (.A(N_809), .B(net_27), .Y(N_69));
    DFN1E1 \scaledatain[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[13]));
    DFN1E1 \noisedata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[4]));
    DFN1E1 \sd_sacq_data[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[6]));
    DFN1E1 \scaleddsdiv[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[0]));
    DFN1E1 dumpload (.D(N_45), .CLK(GLA), .E(net_27), .Q(
        top_code_0_dumpload));
    DFN1E1 \scaledatain[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[7]));
    DFN1E1 \noisedata[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[1]));
    NOR2 n_divnum_1_sqmuxa_0_a2_0_a2 (.A(N_462), .B(N_290), .Y(
        n_divnum_1_sqmuxa));
    DFN1E1 \pd_pluse_data[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[7]));
    DFN1E1 \bri_datain[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[14]));
    DFN1E1 \scandata[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[0]));
    DFN1E1 \n_divnum[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[6]));
    OR2A scanload_3_i_o2_0 (.A(xa_c[7]), .B(un1_xa_7_3), .Y(N_128));
    DFN1E1 \scandata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[6]));
    DFN1E1 \state_1ms_data[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[11]));
    DFN1E1 \scandata[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[1]));
    OR3A un1_state_1ms_rst_n113_2_i_a2_1_o2 (.A(N_268), .B(xa_c[5]), 
        .C(N_278), .Y(N_293));
    DFN1E1 \plusedata[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[1]));
    NOR3 un1_xa_131_2_0_a2_2 (.A(N_232), .B(N_134), .C(xa_c[3]), .Y(
        un1_xa_131_2_0_a2_2_net_1));
    DFN1E1 \sigtimedata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[10]));
    MX2 \relayclose_on_RNO_0[1]  (.A(relayclose_on_c[1]), .B(
        un1_GPMI_0_1_0[1]), .S(relayclose_on_1_sqmuxa), .Y(N_797));
    DFN1E1 \sd_sacq_data[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[9]));
    NOR3B pluse_scale_RNO_5 (.A(N_144_i_0), .B(xa_c[1]), .C(N_134), .Y(
        pluse_scale_3_0_o2_1));
    DFN1 k2 (.D(N_83), .CLK(GLA), .Q(k2_c));
    DFN1E1 \scandata[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[12]));
    OR2A cal_load_3_i_i_o2_0 (.A(xa_c[1]), .B(xa_c[2]), .Y(N_277));
    NOR3A plusedata_1_sqmuxa_0_a2_0_a2 (.A(xa_c_0_7), .B(N_293), .C(
        N_462), .Y(plusedata_1_sqmuxa));
    NOR3 un1_state_1ms_rst_n113_2_i_a2_1_a2 (.A(xa_c_0_7), .B(N_228), 
        .C(N_293), .Y(N_1395));
    DFN1E1 \s_acqnum[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[1]));
    DFN1E1 \dumpdata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[11]));
    DFN1E1 \s_acqnum[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[7]));
    DFN1E1 s_load (.D(N_203), .CLK(GLA), .E(net_27), .Q(
        top_code_0_s_load));
    NOR2 dump_sustain_RNO_2 (.A(N_278), .B(N_282), .Y(
        un1_state_1ms_rst_n113_5_i_a2_0_a2_0));
    NOR3 un1_state_1ms_rst_n113_43_i_a2_2_0 (.A(un1_xa_7_3), .B(
        xa_c[0]), .C(N_233), .Y(N_186_2));
    OR2 dds_choice_3_0_o2_3 (.A(xa_c[2]), .B(xa_c[0]), .Y(N_1559));
    DFN1E1 \noisedata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[7]));
    NOR2 un1_state_1ms_rst_n113_3_i_a2_0_a2 (.A(N_300), .B(N_163_1), 
        .Y(N_163));
    DFN1E1 \pd_pluse_choice[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        pd_pluse_choice_1_sqmuxa), .Q(pd_pluse_choice[2]));
    NOR3 scandata_1_sqmuxa_0_a2_0_a2 (.A(N_288), .B(N_163_1), .C(N_446)
        , .Y(scandata_1_sqmuxa));
    DFN1E1 \state_1ms_data[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[3]));
    DFN1E1 scanchoice (.D(N_12), .CLK(GLA), .E(net_27), .Q(
        top_code_0_scanchoice));
    NOR3C relayclose_on_1_sqmuxa_0_a2_2_a2 (.A(GPMI_0_code_en), .B(
        dumpload_3_i_i_o2_0_net_1), .C(
        relayclose_on_1_sqmuxa_0_a2_2_a2_3_net_1), .Y(
        relayclose_on_1_sqmuxa));
    OR2A scan_start_RNO_3 (.A(N_186_2), .B(N_272), .Y(
        un1_state_1ms_rst_n113_43_i_a2_0));
    AO1A scanload_RNO_1 (.A(N_128), .B(N_159), .C(top_code_0_scanload), 
        .Y(N_194_i));
    DFN1E1 \n_acqnum[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[10]));
    NOR2A un1_state_1ms_rst_n113_28_i_a2_1 (.A(xa_c[4]), .B(N_136), .Y(
        un1_state_1ms_rst_n113_28_i_a2_1_net_1));
    NOR3A change_1_sqmuxa_0_a2_0_a2 (.A(N_459), .B(N_276), .C(N_229), 
        .Y(change_1_sqmuxa));
    OR3B un1_xa_13_0_a2 (.A(N_186_2), .B(xa_c[3]), .C(N_272), .Y(
        un1_xa_13));
    DFN1E1 \sd_sacq_data[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[1]));
    DFN1E1 \state_1ms_lc[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        state_1ms_lc_1_sqmuxa), .Q(state_1ms_lc[1]));
    OR2A n_s_ctrl_3_0_o2_1 (.A(xa_c[0]), .B(N_280), .Y(N_141));
    DFN1E1 \sigtimedata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[6]));
    DFN1E1 \sigtimedata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[4]));
    NOR2B \relayclose_on_RNO[1]  (.A(N_797), .B(net_27), .Y(N_97));
    NOR3B scanchoice_RNO_1 (.A(scanchoice_3_i_a2_0_1), .B(
        scanchoice_3_i_a2_0_0), .C(N_235), .Y(N_197));
    NOR2B pn_change_3_0_o2_0_i_o2 (.A(xa_c[6]), .B(N_269), .Y(N_275));
    DFN1E1 \s_acqnum[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[8]));
    DFN1E1 n_load (.D(N_205), .CLK(GLA), .E(net_27), .Q(
        top_code_0_n_load));
    MX2 \relayclose_on_RNO_0[7]  (.A(relayclose_on_c[7]), .B(
        un1_GPMI_0_1[7]), .S(relayclose_on_1_sqmuxa), .Y(N_803));
    DFN1E1 nstatechoice (.D(N_1543), .CLK(GLA), .E(net_27), .Q(
        top_code_0_nstatechoice));
    DFN1E1 \sigtimedata[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[12]));
    NOR3 scaleload_3_i_i_o2_0 (.A(N_272), .B(N_276), .C(N_229), .Y(
        N_295));
    OAI1 s_load_RNO (.A(N_290), .B(N_296), .C(N_408), .Y(N_203));
    NOR3B dds_choice_RNO_1 (.A(dds_choice_3_0_a2_0_2), .B(
        dds_choice_3_0_a2_0_1), .C(N_140), .Y(N_200));
    OR2A scale_start_RNO_3 (.A(un1_state_1ms_rst_n113_44_i_a2_0_0), .B(
        N_448), .Y(N_351_i));
    DFN1E1 \bri_datain[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[10]));
    NOR3B scale_rst_RNO_3 (.A(xa_c[5]), .B(xa_c[6]), .C(xa_c[2]), .Y(
        un1_state_1ms_rst_n113_35_i_a2_1));
    DFN1E1 bridge_load_0 (.D(N_181), .CLK(GLA), .E(net_27), .Q(
        top_code_0_bridge_load_0));
    AO1 state_1ms_load_RNO_0 (.A(N_160), .B(N_148), .C(
        top_code_0_state_1ms_load), .Y(N_192));
    DFN1E1 sigrst (.D(N_6), .CLK(GLA), .E(net_27), .Q(
        top_code_0_sigrst));
    DFN1E1 \pd_pluse_data[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[14]));
    DFN1E1 \pd_pluse_choice[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        pd_pluse_choice_1_sqmuxa), .Q(pd_pluse_choice[0]));
    OR2B scandata_1_sqmuxa_0_a2_0_a2_0 (.A(xa_c[0]), .B(net_27), .Y(
        N_446));
    DFN1E1 \scandata[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[2]));
    DFN1E1 \plusedata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[10]));
    DFN1E1 \s_addchoice[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        s_addchoice_1_sqmuxa), .Q(s_addchoice[0]));
    NOR2B \relayclose_on_RNO[10]  (.A(N_806), .B(net_27), .Y(N_59));
    MX2A sd_sacq_load_RNO (.A(xa_c[0]), .B(top_code_0_sd_sacq_load), 
        .S(N_310), .Y(N_201));
    DFN1E1 \s_addchoice[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        s_addchoice_1_sqmuxa), .Q(s_addchoice[1]));
    DFN1E1 \n_acqnum[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[11]));
    AO1 noise_start_RNO_2 (.A(un1_state_1ms_rst_n113_43_i_a2_0_1), .B(
        un1_state_1ms_rst_n113_41_i_a2_1), .C(N_123), .Y(
        noise_start_RNO_2_net_1));
    OR2 cal_data_1_sqmuxa_3_0_a2_0_a2 (.A(xa_c[6]), .B(xa_c[5]), .Y(
        un1_xa_7_3));
    NOR3B un1_state_1ms_rst_n113_5_i_a2_0_o2 (.A(GPMI_0_code_en), .B(
        dumpload_3_i_i_o2_0_net_1), .C(xa_c[6]), .Y(N_268));
    OR2A scanload_3_i_o2_1 (.A(xa_c[4]), .B(xa_c[0]), .Y(N_132));
    MX2B scan_start_RNO_0 (.A(top_code_0_scan_start), .B(un1_xa_10), 
        .S(N_31), .Y(N_784));
    OR2A dds_load_3_i_o2_0 (.A(xa_c[0]), .B(N_272), .Y(N_296));
    OR2 scan_start_RNO_5 (.A(N_233), .B(N_277), .Y(
        un1_state_1ms_rst_n113_42_i_a2_1_0));
    OR3C nstatechoice_3_0_i_o2_0 (.A(GPMI_0_code_en), .B(
        nstatechoice_3_0_i_o2_1_m1_e_2_net_1), .C(xa_c[3]), .Y(N_279));
    DFN1E1 \bri_datain[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[3]));
    DFN1E1 \scalechoice[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        scalechoice_1_sqmuxa), .Q(scalechoice[2]));
    DFN1E1 \sigtimedata[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[14]));
    OR3B dumpload_RNO_0 (.A(dumpload_3_i_i_o2_0_net_1), .B(N_156), .C(
        N_158), .Y(N_1562));
    NOR3B halfdata_1_sqmuxa_0_a2_0_a2 (.A(N_287), .B(N_459), .C(N_276), 
        .Y(halfdata_1_sqmuxa));
    DFN1E1 \sd_sacq_data[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[10]));
    DFN1E1 \n_acqnum[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[2]));
    MX2 \relayclose_on_RNO_0[6]  (.A(relayclose_on_c[6]), .B(
        un1_GPMI_0_1[6]), .S(relayclose_on_1_sqmuxa), .Y(N_802));
    DFN1E1 \pd_pluse_data[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[13]));
    DFN1E1 \dumpdata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[8]));
    NOR2A k1_RNO_1 (.A(N_292), .B(N_282), .Y(N_118));
    MX2 \relayclose_on_RNO_0[4]  (.A(relayclose_on_c[4]), .B(
        un1_GPMI_0_1[4]), .S(relayclose_on_1_sqmuxa), .Y(N_800));
    NOR3A noisedata_1_sqmuxa_0_a2_1 (.A(xa_c[4]), .B(N_280), .C(N_122), 
        .Y(noisedata_1_sqmuxa_0_a2_1_net_1));
    OR2A noise_start_RNO_3 (.A(un1_xa_10_0_a2_0_a2_0), .B(N_264), .Y(
        un1_state_1ms_rst_n113_43_i_a2_0_1));
    OR2A change_1_sqmuxa_11_0_a2_0_a2_0_a2_1_a2_0_a2_0 (.A(net_27), .B(
        xa_c_0_0), .Y(N_445));
    NOR3 un1_xa_131_2_0_o2_1 (.A(N_264), .B(N_263), .C(xa_c[11]), .Y(
        N_121));
    NOR2A scanchoice_3_i_o2_1 (.A(xa_c[7]), .B(xa_c[6]), .Y(N_138));
    DFN1E1 \sigtimedata[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[0]));
    NOR2A un1_state_1ms_rst_n113_43_i_a2_11 (.A(N_148), .B(N_122), .Y(
        N_239));
    DFN1 pluse_str (.D(N_87), .CLK(GLA), .Q(top_code_0_pluse_str));
    GND GND_i (.Y(GND));
    NOR2B \relayclose_on_RNO[2]  (.A(N_798), .B(net_27), .Y(N_99));
    NOR2 scale_start_RNO_4 (.A(N_229), .B(xa_c_0_0), .Y(
        un1_state_1ms_rst_n113_44_i_a2_0_0));
    DFN1E1 \state_1ms_data[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[9]));
    DFN1 noise_start (.D(N_85), .CLK(GLA), .Q(top_code_0_noise_start));
    OR2A un1_xa_4_0_o2 (.A(xa_c[2]), .B(xa_c[1]), .Y(N_280));
    DFN1E1 \cal_data[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[4]));
    OR2A un1_state_1ms_rst_n113_3_i_a2_0_a2_1 (.A(xa_c[7]), .B(N_272), 
        .Y(N_163_1));
    OR2B un1_state_1ms_rst_n113_43_i_o2_1 (.A(xa_c[5]), .B(N_125), .Y(
        N_136));
    DFN1E1 \scalechoice[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        scalechoice_1_sqmuxa), .Q(scalechoice[1]));
    DFN1E1 n_s_ctrl_1 (.D(n_s_ctrl_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_n_s_ctrl_1));
    OR2A scaleddsdiv_1_sqmuxa_0_a2_0 (.A(N_287), .B(N_446), .Y(N_451));
    OA1B pluse_noise_ctrl_RNO_0 (.A(N_282), .B(N_300), .C(
        top_code_0_pluse_noise_ctrl), .Y(N_371));
    DFN1E1 \sd_sacq_data[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[7]));
    DFN1E1 \dds_configdata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[9]));
    NOR3B un1_state_1ms_rst_n113_i_a2_0_o2 (.A(N_268), .B(xa_c[5]), .C(
        N_229), .Y(N_292));
    MX2 \relayclose_on_RNO_0[2]  (.A(relayclose_on_c[2]), .B(
        un1_GPMI_0_1_0[2]), .S(relayclose_on_1_sqmuxa), .Y(N_798));
    MX2B noise_start_RNO_0 (.A(top_code_0_noise_start), .B(un1_xa_13), 
        .S(N_29), .Y(N_787));
    NOR3B pd_pluse_choice_1_sqmuxa_0_a2_0_a2 (.A(N_292), .B(xa_c_0_7), 
        .C(N_462), .Y(pd_pluse_choice_1_sqmuxa));
    DFN1E1 dds_choice (.D(dds_choice_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_dds_choice));
    MX2 \relayclose_on_RNO_0[3]  (.A(relayclose_on_c[3]), .B(
        un1_GPMI_0_1[3]), .S(relayclose_on_1_sqmuxa), .Y(N_799));
    DFN1E1 \scandata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[3]));
    DFN1E1 \noisedata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[6]));
    OR2 state_1ms_load_3_i_o2_2 (.A(N_1558), .B(N_122), .Y(N_129));
    DFN1E1 \pd_pluse_data[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[5]));
    DFN1E1 \scalechoice[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        scalechoice_1_sqmuxa), .Q(scalechoice[3]));
    DFN1E1 \scandata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[10]));
    DFN1 \relayclose_on[5]  (.D(N_47), .CLK(GLA), .Q(
        relayclose_on_c[5]));
    NOR2 state_1ms_data_1_sqmuxa_0_a2_0 (.A(N_445), .B(N_228), .Y(
        N_459));
    XOR2 un1_state_1ms_rst_n113_28_i_x2 (.A(xa_c[1]), .B(xa_c[0]), .Y(
        N_120_i));
    DFN1E1 \change_0[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        change_1_sqmuxa), .Q(un1_top_code_0_3_0[0]));
    DFN1E1 \n_divnum[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[5]));
    DFN1 scale_start (.D(N_89), .CLK(GLA), .Q(top_code_0_scale_start));
    DFN1E1 \plusedata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[6]));
    DFN1E1 \plusedata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[11]));
    DFN1E1 \state_1ms_data[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[0]));
    AO1C scaleload_RNO (.A(N_448), .B(scaleload_3_i_i_a2_0_0), .C(
        N_390), .Y(N_175));
    DFN1E1 \pd_pluse_data[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[12]));
    DFN1E1 \cal_data[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[3]));
    DFN1E1 \dumpdata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[7]));
    OR2 n_s_ctrl_3_0_o2_0_0 (.A(N_141), .B(N_147), .Y(
        n_s_ctrl_3_0_o2_0));
    NOR3 s_addchoice_1_sqmuxa_0_a2_0_a2 (.A(N_299), .B(N_228), .C(
        N_458), .Y(s_addchoice_1_sqmuxa));
    DFN1E1 \dds_configdata[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[13]));
    DFN1E1 \scaleddsdiv[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[4]));
    DFN1E1 \n_acqnum[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[3]));
    OA1B dds_load_RNO (.A(N_316), .B(top_code_0_dds_load), .C(N_355), 
        .Y(N_30));
    OR3A state_1ms_start_RNO_2 (.A(xa_c[4]), .B(N_136), .C(N_151), .Y(
        N_190));
    DFN1E1 \dumpdata[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[2]));
    NOR2 sd_sacq_choice_1_sqmuxa_0_a2_0_a2 (.A(
        sd_sacq_choice_1_sqmuxa_1), .B(N_448), .Y(
        sd_sacq_choice_1_sqmuxa));
    AO1C scaleload_RNO_1 (.A(xa_c[0]), .B(N_295), .C(
        top_code_0_scaleload), .Y(N_390));
    OR2A pn_change_RNO_2 (.A(xa_c_0_0), .B(N_278), .Y(
        pn_change_3_0_i_o2_0_net_1));
    DFN1E1 \bri_datain[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[11]));
    OR2 dds_choice_3_0_o2_1 (.A(xa_c[1]), .B(N_123), .Y(N_140));
    OR2A un1_state_1ms_rst_n113_28_i_o2 (.A(GPMI_0_code_en), .B(
        xa_c[3]), .Y(N_1558));
    MX2B k2_RNO_0 (.A(k2_c), .B(xa_c_0_0), .S(N_1449), .Y(N_793));
    DFN1E1 \n_divnum[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[1]));
    DFN1E1 \sigtimedata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[11]));
    NOR2 dds_choice_3_0_o2_0 (.A(xa_c[7]), .B(xa_c[6]), .Y(N_125));
    DFN1E1 \bri_datain[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[9]));
    OR2A un1_xa_30_0_o2 (.A(xa_c[1]), .B(N_1559), .Y(N_158));
    NOR3 un1_xa_49_0_a2 (.A(N_280), .B(N_238), .C(
        un1_xa_49_0_a2_1_net_1), .Y(un1_xa_49));
    DFN1E1 \noisedata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[11]));
    NOR2A scanchoice_RNO_2 (.A(N_138), .B(xa_c[5]), .Y(
        scanchoice_3_i_a2_0_1));
    DFN1 \relayclose_on[15]  (.D(N_73), .CLK(GLA), .Q(
        relayclose_on_c[15]));
    DFN1E1 \scaledatain[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[5]));
    OR2A noise_start_RNO_4 (.A(un1_state_1ms_rst_n113_41_i_a2_1_0), .B(
        N_272), .Y(un1_state_1ms_rst_n113_41_i_a2_1));
    NOR3A pluse_scale_RNO_3 (.A(N_144_i_0), .B(N_262), .C(xa_c[10]), 
        .Y(pluse_scale_3_0_a2_0_0));
    OA1B pd_pluse_load_RNO (.A(N_319), .B(top_code_0_pd_pluse_load), 
        .C(N_395), .Y(N_179));
    NOR3 state_1ms_lc_1_sqmuxa_0_a2_5_a2 (.A(N_299), .B(N_272), .C(
        N_451), .Y(state_1ms_lc_1_sqmuxa));
    DFN1E1 \sigtimedata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[5]));
    DFN1 \relayclose_on[2]  (.D(N_99), .CLK(GLA), .Q(
        relayclose_on_c[2]));
    DFN1E1 \plusedata[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[2]));
    NOR2 scanchoice_RNO_3 (.A(N_122), .B(N_132), .Y(
        scanchoice_3_i_a2_0_0));
    DFN1E1 \sd_sacq_choice[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        sd_sacq_choice_1_sqmuxa), .Q(sd_sacq_choice[3]));
    OR3A dds_choice_RNO_0 (.A(dds_choice_3_0_o2_1_net_1), .B(N_134), 
        .C(N_140), .Y(N_176));
    DFN1E1 \dumpdata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[10]));
    DFN1E1 \n_divnum[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[2]));
    MX2A nstateload_RNO (.A(xa_c[0]), .B(top_code_0_nstateload), .S(
        N_325), .Y(N_82));
    OR2 noisedata_1_sqmuxa_0_o2 (.A(N_128), .B(N_123), .Y(N_157));
    AO1 dds_choice_RNO (.A(top_code_0_dds_choice), .B(N_176), .C(N_200)
        , .Y(dds_choice_3));
    DFN1E1 \scaledatain[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[14]));
    NOR2 pn_change_RNO_1 (.A(pn_change_3_0_i_a2_0_0), .B(N_448), .Y(
        N_393));
    DFN1E1 cal_load (.D(N_106), .CLK(GLA), .E(net_27), .Q(
        top_code_0_cal_load));
    OR2A pn_change_3_0_i_o2_0 (.A(xa_c[3]), .B(xa_c[4]), .Y(N_278));
    DFN1E1 \noisedata[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[0]));
    DFN1E1 \s_acqnum[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[5]));
    DFN1 \relayclose_on[1]  (.D(N_97), .CLK(GLA), .Q(
        relayclose_on_c[1]));
    NOR2A n_load_3_i_i_a2_0_1 (.A(xa_c[0]), .B(N_228), .Y(N_411_1));
    DFN1E1 pluseload (.D(pluseload_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pluseload));
    NOR3B scanload_3_i_o2_2 (.A(xa_c[1]), .B(xa_c[2]), .C(N_129), .Y(
        N_160));
    DFN1E1 \scaledatain[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[8]));
    OR3A nstateload_RNO_0 (.A(xa_c[7]), .B(N_277), .C(N_279), .Y(N_325)
        );
    DFN1E1 \n_acqnum[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[1]));
    NOR2B scan_start_RNO (.A(N_784), .B(net_27), .Y(N_91));
    DFN1E1 \n_acqnum[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[7]));
    NOR3A n_s_ctrl_3_0_a2_0_5 (.A(n_s_ctrl_3_0_a2_0_3_net_1), .B(
        xa_c[16]), .C(xa_c[9]), .Y(n_s_ctrl_3_0_a2_0_5_net_1));
    DFN1E1 \n_divnum[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[9]));
    DFN1E1 bridge_load (.D(N_181), .CLK(GLA), .E(net_27), .Q(
        top_code_0_bridge_load));
    DFN1E1 \cal_data[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[0]));
    DFN1 noise_rst_0_0 (.D(N_38), .CLK(GLA), .Q(top_code_0_noise_rst_0)
        );
    NOR3A un1_xa_2_0_a2 (.A(N_148), .B(N_277), .C(xa_c[3]), .Y(
        un1_xa_2));
    NOR2B pluseload_3_0_o2_1 (.A(N_138), .B(N_130), .Y(N_144_i_0));
    NOR2 acqclken_3_0_o2_0_0 (.A(acqclken_3_0_o2_0_0_1_net_1), .B(
        acqclken_3_0_o2_0_0_0_net_1), .Y(N_260));
    OR2A state_1ms_rst_n_RNIP6MA3 (.A(net_27), .B(N_788), .Y(N_225));
    AO1B scale_start_RNO_1 (.A(N_327), .B(GPMI_0_code_en), .C(N_351_i), 
        .Y(N_26));
    DFN1E1 \change[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        change_1_sqmuxa), .Q(change[0]));
    DFN1 \relayclose_on[11]  (.D(N_62), .CLK(GLA), .Q(
        relayclose_on_c[11]));
    DFN1 \relayclose_on[14]  (.D(N_71), .CLK(GLA), .Q(
        relayclose_on_c[14]));
    DFN1E1 acqclken (.D(acqclken_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_acqclken));
    DFN1E1 \s_addchoice[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        s_addchoice_1_sqmuxa), .Q(s_addchoice[3]));
    DFN1E1 \s_acqnum[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[13]));
    OR2A sigtimedata_1_sqmuxa_0_o2 (.A(xa_c[7]), .B(N_228), .Y(N_282));
    DFN1E1 \scandata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[7]));
    DFN1 \relayclose_on[7]  (.D(N_52), .CLK(GLA), .Q(
        relayclose_on_c[7]));
    DFN1E1 \dumpdata[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[0]));
    DFN1E1 \sigtimedata[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[13]));
    DFN1E1 \sigtimedata[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[1]));
    DFN1E1 \state_1ms_data[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[15]));
    NOR2B \relayclose_on_RNO[12]  (.A(N_808), .B(net_27), .Y(N_66));
    DFN1E1 \n_acqnum[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[8]));
    DFN1E1 \noisedata[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[2]));
    DFN1E1 \scalechoice[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        scalechoice_1_sqmuxa), .Q(scalechoice[4]));
    OR3C state_1ms_start_RNO_1 (.A(N_191), .B(N_352), .C(N_190), .Y(
        N_1554));
    DFN1E1 \state_1ms_data[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[10]));
    OR2A acqclken_3_0_o2_0 (.A(xa_c[4]), .B(N_141), .Y(N_150));
    DFN1E1 \scandata[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[13]));
    DFN1 pluse_rst (.D(N_41), .CLK(GLA), .Q(top_code_0_pluse_rst));
    OR3A sd_sacq_load_RNO_0 (.A(N_287), .B(N_272), .C(N_276), .Y(N_310)
        );
    DFN1E1 \bri_datain[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[1]));
    DFN1E1 \cal_data[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[2]));
    NOR2B \relayclose_on_RNO[11]  (.A(N_807), .B(net_27), .Y(N_62));
    DFN1 state_1ms_rst_n (.D(N_225), .CLK(GLA), .Q(
        top_code_0_state_1ms_rst_n));
    DFN1E1 \sd_sacq_data[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[2]));
    DFN1E1 state_1ms_load (.D(state_1ms_load_RNO_net_1), .CLK(GLA), .E(
        net_27), .Q(top_code_0_state_1ms_load));
    NOR3 n_s_ctrl_3_0_a2_0_0 (.A(N_262), .B(xa_c[10]), .C(N_232), .Y(
        n_s_ctrl_3_0_a2_0_0_net_1));
    DFN1E1 \s_periodnum[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        s_periodnum_1_sqmuxa), .Q(s_periodnum[2]));
    OR3C noise_start_RNO_1 (.A(N_188), .B(noise_start_RNO_2_net_1), .C(
        N_31_2), .Y(N_29));
    NOR2 pluseload_3_0_o2_2 (.A(xa_c[5]), .B(xa_c[4]), .Y(N_130));
    MX2 \relayclose_on_RNO_0[11]  (.A(relayclose_on_c[11]), .B(
        un1_GPMI_0_1[11]), .S(relayclose_on_1_sqmuxa), .Y(N_807));
    NOR3B acqclken_RNO_3 (.A(N_121), .B(acqclken_3_0_o2_1), .C(N_132), 
        .Y(acqclken_3_0_o2_2));
    NOR2A scaleload_RNO_0 (.A(xa_c_0_0), .B(N_229), .Y(
        scaleload_3_i_i_a2_0_0));
    NOR2 n_rd_en_RNO_1 (.A(N_297), .B(N_290), .Y(N_386));
    DFN1 state_1ms_rst_n_0_0 (.D(N_225), .CLK(GLA), .Q(
        top_code_0_state_1ms_rst_n_0));
    DFN1E1 \sigtimedata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[3]));
    OR2 dump_cho_1_sqmuxa_2_0_a2_0_o2_i_a2 (.A(xa_c[2]), .B(xa_c[1]), 
        .Y(N_228));
    NOR2 scale_rst_RNO_1 (.A(xa_c[3]), .B(N_158), .Y(un1_xa_30));
    MX2B k1_RNO_0 (.A(k1_c), .B(xa_c_0_0), .S(N_118), .Y(N_794));
    DFN1E1 \pd_pluse_data[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[15]));
    DFN1E1 n_s_ctrl (.D(n_s_ctrl_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_n_s_ctrl));
    NOR3 bri_datain_1_sqmuxa_0_a2_0_a2 (.A(N_272), .B(N_276), .C(N_458)
        , .Y(bri_datain_1_sqmuxa));
    DFN1E1 \sd_sacq_data[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[14]));
    DFN1E1 \pd_pluse_data[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[2]));
    DFN1E1 \bri_datain[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[4]));
    MX2 \relayclose_on_RNO_0[9]  (.A(relayclose_on_c[9]), .B(
        un1_GPMI_0_1[9]), .S(relayclose_on_1_sqmuxa), .Y(N_805));
    NOR2A pn_change_3_0_o2_0_i_o2_0 (.A(xa_c[5]), .B(xa_c[7]), .Y(
        N_269));
    OR2 un1_state_1ms_rst_n113_43_i_a2_6 (.A(N_232), .B(N_122), .Y(
        N_233));
    OA1 un1_state_1ms_rst_n113_41_i_2 (.A(N_151), .B(
        un1_state_1ms_rst_n113_43_i_a2_2_0_net_1), .C(N_191), .Y(
        N_31_2));
    DFN1E1 \state_1ms_data[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[5]));
    OR2 un1_state_1ms_rst_n113_44_i_a2_1 (.A(N_280), .B(N_276), .Y(
        N_448));
    DFN1E1 \halfdata[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[2]));
    NOR3 n_acqnum_1_sqmuxa_0_a2_0_a2 (.A(N_446), .B(N_277), .C(N_290), 
        .Y(n_acqnum_1_sqmuxa));
    NOR3 dump_cho_1_sqmuxa_0_a2_0_a2 (.A(N_276), .B(N_228), .C(N_451), 
        .Y(dump_cho_1_sqmuxa));
    DFN1E1 \bri_datain[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[15]));
    OAI1 s_load_RNO_0 (.A(N_299), .B(N_309), .C(top_code_0_s_load), .Y(
        N_408));
    DFN1E1 \noisedata[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[14]));
    DFN1E1 \plusedata[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[15]));
    OR3B sigrst_3_i_o2_0 (.A(GPMI_0_code_en), .B(
        nstatechoice_3_0_i_o2_1_m1_e_2_net_1), .C(xa_c[3]), .Y(N_288));
    NOR2B un1_xa_131_3_1 (.A(un1_xa_10), .B(un1_xa_13), .Y(
        un1_xa_131_3_1_net_1));
    AO1A acqclken_RNO (.A(N_123), .B(acqclken_3_0_a2_0_3), .C(N_219), 
        .Y(acqclken_3));
    NOR3 dds_load_RNO_1 (.A(N_288), .B(xa_c_0_7), .C(N_296), .Y(N_355));
    DFN1E1 \sd_sacq_choice[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        sd_sacq_choice_1_sqmuxa), .Q(sd_sacq_choice[1]));
    DFN1E1 \s_acqnum[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[11]));
    OR3B scale_start_RNO_2 (.A(un1_xa_131_3_0_net_1), .B(
        un1_xa_131_3_1_net_1), .C(un1_xa_49), .Y(N_327));
    DFN1E1 \scaleddsdiv[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[3]));
    DFN1E1 \dds_configdata[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[2]));
    OR2 un1_state_1ms_rst_n113_43_i_a2_8 (.A(N_1558), .B(N_280), .Y(
        N_235));
    DFN1E1 \pd_pluse_data[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[10]));
    NOR2B k2_RNO (.A(N_793), .B(net_27), .Y(N_83));
    NOR2B k1_RNO (.A(N_794), .B(net_27), .Y(N_81));
    OA1B sigrst_RNO (.A(N_317), .B(top_code_0_sigrst), .C(N_341), .Y(
        N_6));
    DFN1E1 \s_acqnum[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[15]));
    NOR3A noisedata_1_sqmuxa_0_a2 (.A(noisedata_1_sqmuxa_0_a2_1_net_1), 
        .B(N_157), .C(N_445), .Y(noisedata_1_sqmuxa));
    DFN1E1 \dumpdata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[3]));
    DFN1E1 \plusedata[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[14]));
    DFN1E1 \n_divnum[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[8]));
    DFN1E1 scanload (.D(N_1556_i_0), .CLK(GLA), .E(net_27), .Q(
        top_code_0_scanload));
    OR3B dumpload_RNO_1 (.A(N_411_1), .B(N_156), .C(N_122), .Y(N_222));
    OA1A pluse_scale_RNO_1 (.A(pluse_scale_3_0_o2_1), .B(N_1558), .C(
        top_code_0_pluse_scale), .Y(N_215));
    DFN1E1 n_s_ctrl_0 (.D(n_s_ctrl_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_n_s_ctrl_0));
    DFN1E1 \n_divnum[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[4]));
    NOR2B \relayclose_on_RNO[9]  (.A(N_805), .B(net_27), .Y(N_56));
    NOR2B state_1ms_start_RNO (.A(N_783), .B(net_27), .Y(N_93));
    DFN1E1 \scaledatain[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[12]));
    DFN1E1 \pd_pluse_data[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[6]));
    DFN1E1 \scaledatain[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[15]));
    DFN1E1 \pd_pluse_data[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[1]));
    DFN1E1 \s_acqnum[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[9]));
    DFN1E1 \s_acqnum[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[0]));
    AO1C n_load_RNO (.A(N_290), .B(N_411_1), .C(N_410), .Y(N_205));
    DFN1E1 \s_acqnum[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[14]));
    DFN1E1 \dumpdata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[4]));
    NOR2 n_rd_en_RNO_0 (.A(N_296), .B(N_286), .Y(N_320));
    DFN1E1 \dumpdata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[5]));
    DFN1E1 \dds_configdata[14]  (.D(un1_GPMI_0_1[14]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[14]));
    DFN1E1 \scaledatain[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[2]));
    DFN1E1 \s_acqnum[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[4]));
    DFN1E1 \bri_datain[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[6]));
    DFN1E1 \plusedata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[9]));
    DFN1E1 \dump_cho[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        dump_cho_1_sqmuxa), .Q(dump_cho[1]));
    DFN1E1 \halfdata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[6]));
    DFN1E1 \dds_configdata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[11]));
    OR2 acqclken_3_0_o2_0_0_1 (.A(xa_c[14]), .B(xa_c[15]), .Y(
        acqclken_3_0_o2_0_0_1_net_1));
    DFN1E1 \pd_pluse_data[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[4]));
    OA1B RAM_Rd_rst_RNO_0 (.A(N_272), .B(N_294), .C(
        top_code_0_RAM_Rd_rst), .Y(N_381));
    AO1C pluseload_RNO (.A(N_1565), .B(top_code_0_pluseload), .C(N_214)
        , .Y(pluseload_3));
    OR2 pd_pluse_choice_1_sqmuxa_0_a2_0_a2_0 (.A(N_445), .B(N_280), .Y(
        N_462));
    DFN1E1 \scaledatain[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[10]));
    DFN1 noise_rst (.D(N_38), .CLK(GLA), .Q(top_code_0_noise_rst));
    NOR2 nstatechoice_3_0_i_o2_1_m1_e_1 (.A(xa_c[5]), .B(xa_c[6]), .Y(
        nstatechoice_3_0_i_o2_1_m1_e_1_net_1));
    MX2 \relayclose_on_RNO_0[8]  (.A(relayclose_on_c[8]), .B(
        un1_GPMI_0_1[8]), .S(relayclose_on_1_sqmuxa), .Y(N_804));
    OR2A un1_state_1ms_rst_n113_43_i_a2_1 (.A(N_239), .B(N_235), .Y(
        N_188));
    NOR2B \relayclose_on_RNO[8]  (.A(N_804), .B(net_27), .Y(N_54));
    DFN1E1 \halfdata[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[1]));
    DFN1E1 \pd_pluse_choice[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        pd_pluse_choice_1_sqmuxa), .Q(pd_pluse_choice[3]));
    MX2 pluse_str_RNO_0 (.A(top_code_0_pluse_str), .B(un1_xa_49), .S(
        N_28), .Y(N_786));
    NOR3 relayclose_on_1_sqmuxa_0_a2_2_a2_2 (.A(N_297), .B(N_229), .C(
        xa_c_0_7), .Y(relayclose_on_1_sqmuxa_0_a2_2_a2_2_net_1));
    NOR2A pluse_str_RNO_2 (.A(xa_c_0_7), .B(N_280), .Y(
        un1_state_1ms_rst_n113_45_i_a2_0_0));
    DFN1E1 \noisedata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[5]));
    NOR2A sigrst_RNO_0 (.A(N_303), .B(N_288), .Y(N_317));
    OR3C scan_start_RNO_1 (.A(N_188), .B(un1_state_1ms_rst_n113_42_i_0)
        , .C(N_31_2), .Y(N_31));
    NOR3C pluse_scale_RNO_0 (.A(pluse_scale_3_0_a2_0_1), .B(
        pluse_scale_3_0_a2_0_0), .C(pluse_scale_3_0_a2_0_2), .Y(
        pluse_scale_3_0_a2_0_4));
    MX2 scan_rst_0_0_RNICPJQ2 (.A(net_33_0), .B(xa_c_0_0), .S(N_1395), 
        .Y(N_790));
    DFN1E1 \state_1ms_data[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[13]));
    NOR2 dumpload_3_i_i_o2_0_1 (.A(N_264), .B(N_220_1_i_0), .Y(
        dumpload_3_i_i_o2_0_net_1));
    NOR3 un1_state_1ms_rst_n113_1_i_a2_0_a2 (.A(xa_c_0_7), .B(N_280), 
        .C(N_293), .Y(N_164));
    DFN1 \relayclose_on[10]  (.D(N_59), .CLK(GLA), .Q(
        relayclose_on_c[10]));
    OR2B scalechoice_1_sqmuxa_0_a2_2_i_o2 (.A(xa_c[2]), .B(xa_c[1]), 
        .Y(N_272));
    OR3A un1_state_1ms_rst_n113_45_i_o2_0 (.A(N_268), .B(xa_c[5]), .C(
        N_229), .Y(N_300));
    NOR3 s_periodnum_1_sqmuxa_0_a2_0_a2 (.A(N_445), .B(N_272), .C(
        N_290), .Y(s_periodnum_1_sqmuxa));
    DFN1E1 \noisedata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[9]));
    DFN1E1 \state_1ms_data[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[4]));
    DFN1 scale_rst (.D(N_223), .CLK(GLA), .Q(scale_rst_net_1));
    OR2A noise_rst_0_0_RNID5DS2 (.A(net_27), .B(N_792), .Y(N_38));
    DFN1E1 \sd_sacq_data[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[12]));
    DFN1E1 \scandata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[4]));
    DFN1E1 \scaleddsdiv[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[1]));
    MX2B dump_sustain_RNO_0 (.A(top_code_0_dump_sustain), .B(xa_c_0_0), 
        .S(N_119), .Y(N_795));
    DFN1E1 dds_load (.D(N_30), .CLK(GLA), .E(net_27), .Q(
        dds_load_net_1));
    DFN1E1 \scaledatain[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[11]));
    NOR2 n_s_ctrl_3_0_a2_0_3 (.A(xa_c[17]), .B(xa_c[18]), .Y(
        n_s_ctrl_3_0_a2_0_3_net_1));
    NOR3 n_s_ctrl_3_0_a2_0_1 (.A(un1_xa_7_3), .B(xa_c_0_0), .C(xa_c[8])
        , .Y(n_s_ctrl_3_0_a2_0_1_net_1));
    DFN1E1 \state_1ms_data[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[2]));
    AO1B dumpload_RNO (.A(top_code_0_dumpload), .B(N_1562), .C(N_222), 
        .Y(N_45));
    DFN1E1 \scalechoice[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        scalechoice_1_sqmuxa), .Q(scalechoice[0]));
    NOR3C nstatechoice_3_0_i_o2_1_m1_e_2 (.A(xa_c[4]), .B(
        dumpload_3_i_i_o2_0_net_1), .C(
        nstatechoice_3_0_i_o2_1_m1_e_1_net_1), .Y(
        nstatechoice_3_0_i_o2_1_m1_e_2_net_1));
    CLKINT scale_rst_RNIA6G4 (.A(scale_rst_net_1), .Y(
        top_code_0_scale_rst));
    NOR3B dumpload_3_i_i_o2_0 (.A(N_275), .B(GPMI_0_code_en), .C(N_278)
        , .Y(N_156));
    OR3B un1_state_1ms_rst_n113_43_i_a2_2_0_0 (.A(xa_c[5]), .B(xa_c[6])
        , .C(N_232), .Y(un1_state_1ms_rst_n113_43_i_a2_2_0_net_1));
    DFN1E1 \state_1ms_lc[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        state_1ms_lc_1_sqmuxa), .Q(state_1ms_lc[3]));
    DFN1E1 nstateload (.D(N_82), .CLK(GLA), .E(net_27), .Q(
        top_code_0_nstateload));
    NOR2A dds_choice_RNO_4 (.A(xa_c[4]), .B(N_1559), .Y(
        dds_choice_3_0_a2_0_1));
    DFN1E1 \sd_sacq_data[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[3]));
    OR2 bridge_load_3_0_i_o2_1 (.A(N_297), .B(N_278), .Y(N_309));
    OR3A un1_state_1ms_rst_n113_43_i_o2_3 (.A(xa_c[1]), .B(N_129), .C(
        N_124), .Y(N_151));
    DFN1E1 \state_1ms_lc[0]  (.D(un1_GPMI_0_1[0]), .CLK(GLA), .E(
        state_1ms_lc_1_sqmuxa), .Q(state_1ms_lc[0]));
    NOR3 scalechoice_1_sqmuxa_0_a2_0_a2 (.A(N_272), .B(N_276), .C(
        scalechoice_1_sqmuxa_0_a2_0_a2_0_net_1), .Y(
        scalechoice_1_sqmuxa));
    DFN1E1 \scandata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[9]));
    DFN1E1 \dds_configdata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[3]));
    DFN1E1 pluse_lc (.D(N_70), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pluse_lc));
    OR3 un1_state_1ms_rst_n113_43_i_a2_4 (.A(xa_c_0_0), .B(N_238), .C(
        N_235), .Y(N_191));
    DFN1E1 \pd_pluse_data[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[11]));
    DFN1E1 \n_acqnum[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[5]));
    DFN1E1 \state_1ms_data[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[7]));
    DFN1E1 \pd_pluse_data[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[0]));
    NOR2 sigrst_RNO_1 (.A(sigrst_3_i_a2_0_0), .B(N_288), .Y(N_341));
    OA1B pn_change_RNO (.A(N_315), .B(top_code_0_pn_change), .C(N_393), 
        .Y(N_177));
    NOR3B k2_RNO_1 (.A(xa_c_0_7), .B(N_292), .C(N_277), .Y(N_1449));
    DFN1E1 \dump_cho[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        dump_cho_1_sqmuxa), .Q(dump_cho[2]));
    DFN1E1 \change_0[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        change_1_sqmuxa), .Q(un1_top_code_0_3_0[1]));
    DFN1E1 \sigtimedata[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[15]));
    DFN1E1 \halfdata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[3]));
    OR2B state_1ms_data_1_sqmuxa_0_o2 (.A(N_269), .B(N_268), .Y(N_299));
    DFN1E1 \sd_sacq_data[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[13]));
    OA1B nstatechoice_RNO_0 (.A(N_279), .B(N_282), .C(
        top_code_0_nstatechoice), .Y(N_377));
    DFN1 k1 (.D(N_81), .CLK(GLA), .Q(k1_c));
    DFN1E1 \plusedata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[5]));
    OR2 un1_state_1ms_rst_n113_2_0_i_0_a2_0_a2_0_o2_i_a2 (.A(xa_c[4]), 
        .B(xa_c[3]), .Y(N_229));
    MX2 \relayclose_on_RNO_0[12]  (.A(relayclose_on_c[12]), .B(
        un1_GPMI_0_1[12]), .S(relayclose_on_1_sqmuxa), .Y(N_808));
    DFN1 pluse_rst_0_0 (.D(N_41), .CLK(GLA), .Q(top_code_0_pluse_rst_0)
        );
    NOR2B \relayclose_on_RNO[5]  (.A(N_801), .B(net_27), .Y(N_47));
    AOI1B un1_xa_131_3_0 (.A(un1_xa_131_2_0_a2_2_net_1), .B(
        un1_xa_131_2_0_a2_1_net_1), .C(un1_xa_4), .Y(
        un1_xa_131_3_0_net_1));
    OR3A un1_xa_4_0_a2 (.A(N_239), .B(N_280), .C(xa_c[3]), .Y(un1_xa_4)
        );
    OR2A scale_rst_RNO (.A(net_27), .B(N_789), .Y(N_223));
    NOR2A scale_rst_RNO_4 (.A(N_120_i), .B(N_233), .Y(
        un1_state_1ms_rst_n113_35_i_a2_0));
    DFN1E1 \pd_pluse_choice[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        pd_pluse_choice_1_sqmuxa), .Q(pd_pluse_choice[1]));
    NOR3C dump_sustain_RNO_1 (.A(un1_state_1ms_rst_n113_5_i_a2_0_a2_0), 
        .B(xa_c[5]), .C(N_268), .Y(N_119));
    DFN1E1 \dds_configdata[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[6]));
    NOR3A acqclken_RNO_2 (.A(N_138), .B(N_150), .C(xa_c[5]), .Y(
        acqclken_3_0_a2_0_2));
    OR2 pluseload_3_0_o2_3 (.A(N_124), .B(N_122), .Y(N_134));
    OA1B RAM_Rd_rst_RNO (.A(N_141), .B(N_286), .C(N_381), .Y(N_1544));
    DFN1 \relayclose_on[6]  (.D(N_50), .CLK(GLA), .Q(
        relayclose_on_c[6]));
    DFN1E1 \sd_sacq_data[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[8]));
    DFN1E1 \sd_sacq_choice[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        sd_sacq_choice_1_sqmuxa), .Q(sd_sacq_choice[2]));
    DFN1E1 \state_1ms_data[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[12]));
    NOR2A acqclken_RNO_4 (.A(N_260), .B(N_272), .Y(acqclken_3_0_o2_1));
    OR2 acqclken_3_0_o2_0_0_0 (.A(xa_c[12]), .B(xa_c[13]), .Y(
        acqclken_3_0_o2_0_0_0_net_1));
    OR2 cal_load_3_i_i_o2_2 (.A(xa_c[0]), .B(N_286), .Y(N_294));
    NOR3 un1_state_1ms_rst_n113_43_i_a2_0_1_0_0 (.A(N_158), .B(
        N_220_1_i_0), .C(N_147), .Y(un1_xa_10_0_a2_0_a2_0));
    DFN1E1 \scaleddsdiv[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[2]));
    NOR3B un1_state_1ms_rst_n113_28_i_a2 (.A(
        un1_state_1ms_rst_n113_28_i_a2_2_net_1), .B(
        un1_state_1ms_rst_n113_28_i_a2_1_net_1), .C(N_1558), .Y(N_209));
    OR2A un1_state_1ms_rst_n113_43_i_a2_10 (.A(N_144_i_0), .B(N_122), 
        .Y(N_238));
    OA1A acqclken_RNO_1 (.A(acqclken_3_0_o2_2), .B(N_157), .C(
        top_code_0_acqclken), .Y(N_219));
    NOR3A un1_state_1ms_rst_n113_28_i_a2_2 (.A(N_120_i), .B(N_122), .C(
        xa_c[2]), .Y(un1_state_1ms_rst_n113_28_i_a2_2_net_1));
    OR3 un1_xa_48_11_0_a2_0_a2_0_o2 (.A(xa_c[9]), .B(xa_c[8]), .C(
        xa_c[10]), .Y(N_263));
    DFN1E1 \n_divnum[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[3]));
    DFN1E1 \noisedata[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[15]));
    AOI1 bridge_load_0_RNIAKBO2 (.A(xa_c_0_0), .B(N_295), .C(
        top_code_0_bridge_load_0), .Y(N_396));
    OA1C nstatechoice_RNO (.A(N_303), .B(N_279), .C(N_377), .Y(N_1543));
    OR2 pn_change_RNO_3 (.A(N_278), .B(xa_c_0_0), .Y(
        pn_change_3_0_i_a2_0_0));
    NOR3 scaleddsdiv_1_sqmuxa_0_a2 (.A(N_276), .B(N_277), .C(N_451), 
        .Y(scaleddsdiv_1_sqmuxa));
    DFN1E1 \plusedata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[4]));
    OR2 n_rd_en_3_0_i_o2_1 (.A(xa_c[0]), .B(N_228), .Y(N_297));
    OR2B un1_state_1ms_rst_n113_43_i_o2_2 (.A(N_130), .B(N_125), .Y(
        N_147));
    DFN1E1 \scaledatain[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[1]));
    DFN1E1 \halfdata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[5]));
    NOR2B \relayclose_on_RNO[3]  (.A(N_799), .B(net_27), .Y(N_101));
    GND GND_i_0 (.Y(GND_0));
    NOR2 scaledatain_1_sqmuxa_0_a2_0_a2 (.A(N_458), .B(N_448), .Y(
        scaledatain_1_sqmuxa));
    DFN1E1 \n_divnum[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        n_divnum_1_sqmuxa), .Q(n_divnum[0]));
    DFN1 \relayclose_on[12]  (.D(N_66), .CLK(GLA), .Q(
        relayclose_on_c[12]));
    AO1B un1_state_1ms_rst_n113_45_i_a2 (.A(un1_xa_131_3_1_net_1), .B(
        un1_xa_131_3_0_net_1), .C(GPMI_0_code_en), .Y(N_352));
    DFN1E1 \scaledatain[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[9]));
    NOR3 pn_change_RNO_0 (.A(N_276), .B(N_277), .C(
        pn_change_3_0_i_o2_0_net_1), .Y(N_315));
    MX2 \relayclose_on_RNO_0[15]  (.A(relayclose_on_c[15]), .B(
        un1_GPMI_0_1[15]), .S(relayclose_on_1_sqmuxa), .Y(N_811));
    NOR2A s_acqnum_1_sqmuxa_0_a2_0_a2 (.A(N_461), .B(N_290), .Y(
        s_acqnum_1_sqmuxa));
    DFN1 scan_rst (.D(N_43), .CLK(GLA), .Q(net_33));
    DFN1E1 \s_acqnum[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[6]));
    DFN1E1 \noisedata[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[3]));
    NOR3C n_s_ctrl_3_0_a2_0_6 (.A(n_s_ctrl_3_0_a2_0_1_net_1), .B(
        n_s_ctrl_3_0_a2_0_0_net_1), .C(n_s_ctrl_3_0_a2_0_5_net_1), .Y(
        n_s_ctrl_3_0_a2_0_6_net_1));
    MX2 scale_rst_RNO_0 (.A(top_code_0_scale_rst), .B(un1_xa_30), .S(
        N_210), .Y(N_789));
    DFN1E1 \scandata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[8]));
    MX2 \relayclose_on_RNO_0[14]  (.A(relayclose_on_c[14]), .B(
        un1_GPMI_0_1[14]), .S(relayclose_on_1_sqmuxa), .Y(N_810));
    DFN1E1 \bri_datain[2]  (.D(un1_GPMI_0_1_0[2]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[2]));
    NOR3A dds_choice_RNO_3 (.A(N_125), .B(N_122), .C(xa_c[5]), .Y(
        dds_choice_3_0_a2_0_2));
    NOR3B pd_pluse_load_RNO_1 (.A(N_292), .B(xa_c_0_7), .C(N_296), .Y(
        N_395));
    OR2 acqclken_3_0_a2_0_1 (.A(N_263), .B(N_262), .Y(N_220_1_i_0));
    DFN1E1 \scandata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[5]));
    DFN1E1 \dds_configdata[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[1]));
    DFN1E1 \dumpdata[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[1]));
    OR2B un1_state_1ms_rst_n113_43_i_o2 (.A(xa_c[3]), .B(
        GPMI_0_code_en), .Y(N_123));
    DFN1E1 \bri_datain[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[13]));
    OR2 scanload_RNO_0 (.A(N_128), .B(N_132), .Y(scanload_3_i_a2_0_0));
    DFN1E1 \plusedata[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        plusedata_1_sqmuxa), .Q(plusedata[12]));
    NOR2 noise_start_RNO_5 (.A(N_122), .B(N_147), .Y(
        un1_state_1ms_rst_n113_41_i_a2_1_0));
    NOR3B state_1ms_data_1_sqmuxa_0_a2 (.A(
        state_1ms_data_1_sqmuxa_0_a2_0_net_1), .B(N_459), .C(N_299), 
        .Y(state_1ms_data_1_sqmuxa));
    DFN1E1 \change[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        change_1_sqmuxa), .Q(change[1]));
    DFN1E1 \n_acqnum[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[9]));
    DFN1E1 \n_acqnum[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[0]));
    DFN1E1 \halfdata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[4]));
    DFN1E1 \state_1ms_data[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[1]));
    OR3 un1_state_1ms_rst_n113_43_i_o2_0 (.A(xa_c[17]), .B(xa_c[16]), 
        .C(xa_c[18]), .Y(N_264));
    DFN1E1 n_rd_en (.D(N_168), .CLK(GLA), .E(net_27), .Q(
        top_code_0_n_rd_en));
    DFN1E1 \n_acqnum[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        n_acqnum_1_sqmuxa), .Q(n_acqnum[4]));
    NOR3 sigtimedata_1_sqmuxa_0_a2 (.A(N_288), .B(N_282), .C(N_445), 
        .Y(sigtimedata_1_sqmuxa));
    DFN1E1 \bri_datain[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[8]));
    OR2A scan_rst_0_0_RNI47ES2 (.A(net_27), .B(N_790), .Y(N_43));
    NOR3B relayclose_on_1_sqmuxa_0_a2_2_a2_3 (.A(xa_c[6]), .B(
        relayclose_on_1_sqmuxa_0_a2_2_a2_2_net_1), .C(xa_c[5]), .Y(
        relayclose_on_1_sqmuxa_0_a2_2_a2_3_net_1));
    MX2 state_1ms_rst_n_RNI1PR83 (.A(top_code_0_state_1ms_rst_n), .B(
        un1_xa_2), .S(N_209), .Y(N_788));
    NOR2 pluse_scale_RNO_2 (.A(N_158), .B(N_264), .Y(
        pluse_scale_3_0_a2_0_1));
    DFN1 \relayclose_on[3]  (.D(N_101), .CLK(GLA), .Q(
        relayclose_on_c[3]));
    DFN1E1 \cal_data[1]  (.D(un1_GPMI_0_1_0[1]), .CLK(GLA), .E(
        cal_data_1_sqmuxa), .Q(cal_data[1]));
    DFN1 scan_rst_0_0 (.D(N_43), .CLK(GLA), .Q(net_33_0));
    NOR3 dds_load_RNO_0 (.A(N_288), .B(xa_c[7]), .C(N_272), .Y(N_316));
    NOR2B \relayclose_on_RNO[14]  (.A(N_810), .B(net_27), .Y(N_71));
    NOR3A dds_choice_RNO_2 (.A(xa_c[4]), .B(xa_c_0_7), .C(un1_xa_7_3), 
        .Y(dds_choice_3_0_o2_1_net_1));
    DFN1E1 \dumpdata[9]  (.D(un1_GPMI_0_1[9]), .CLK(GLA), .E(
        dumpdata_1_sqmuxa), .Q(dumpdata[9]));
    DFN1 scan_start (.D(N_91), .CLK(GLA), .Q(top_code_0_scan_start));
    NOR3C pd_pluse_data_1_sqmuxa_0_a2_0_a2 (.A(N_292), .B(xa_c_0_7), 
        .C(N_461), .Y(pd_pluse_data_1_sqmuxa));
    DFN1E1 \state_1ms_lc[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        state_1ms_lc_1_sqmuxa), .Q(state_1ms_lc[2]));
    DFN1E1 \dds_configdata[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[10]));
    NOR3C un1_xa_131_2_0_a2_1 (.A(xa_c[5]), .B(xa_c[6]), .C(xa_c[1]), 
        .Y(un1_xa_131_2_0_a2_1_net_1));
    NOR2B \relayclose_on_RNO[6]  (.A(N_802), .B(net_27), .Y(N_50));
    DFN1E1 \dump_cho[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        dump_cho_1_sqmuxa), .Q(dump_cho[0]));
    DFN1E1 \noisedata[13]  (.D(un1_GPMI_0_1[13]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[13]));
    DFN1E1 pn_change (.D(N_177), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pn_change));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 dump_sustain (.D(N_79), .CLK(GLA), .Q(top_code_0_dump_sustain)
        );
    DFN1E1 scaleload (.D(N_175), .CLK(GLA), .E(net_27), .Q(
        top_code_0_scaleload));
    NOR2 state_1ms_load_3_i_o2_1 (.A(N_150), .B(N_129), .Y(N_159));
    OR3C bridge_load_3_0_i_o2_0 (.A(GPMI_0_code_en), .B(
        dumpload_3_i_i_o2_0_net_1), .C(N_275), .Y(N_276));
    AO1C pluse_str_RNO_1 (.A(N_300), .B(
        un1_state_1ms_rst_n113_45_i_a2_0_0), .C(N_352), .Y(N_28));
    DFN1E1 \s_periodnum[1]  (.D(un1_GPMI_0_1[1]), .CLK(GLA), .E(
        s_periodnum_1_sqmuxa), .Q(s_periodnum[1]));
    OR2A pluse_rst_RNIEHKS2 (.A(net_27), .B(N_791), .Y(N_41));
    DFN1E1 \dds_configdata[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[5]));
    NOR2B scale_start_RNO (.A(N_785), .B(net_27), .Y(N_89));
    NOR3A acqclken_RNO_0 (.A(acqclken_3_0_a2_0_2), .B(N_264), .C(
        N_220_1_i_0), .Y(acqclken_3_0_a2_0_3));
    DFN1E1 \bri_datain[0]  (.D(un1_GPMI_0_1_0[0]), .CLK(GLA), .E(
        bri_datain_1_sqmuxa), .Q(bri_datain[0]));
    NOR3A dds_configdata_1_sqmuxa_0_a2_0_a2 (.A(N_461), .B(N_288), .C(
        xa_c[7]), .Y(dds_configdata_1_sqmuxa));
    DFN1 \relayclose_on[8]  (.D(N_54), .CLK(GLA), .Q(
        relayclose_on_c[8]));
    DFN1E1 \sd_sacq_data[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[15]));
    DFN1E1 \dds_configdata[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[12]));
    DFN1E1 \state_1ms_data[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[8]));
    NOR2A pluse_noise_ctrl_3_0_i_o2_0 (.A(xa_c[0]), .B(N_282), .Y(
        N_303));
    DFN1E1 \scandata[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        scandata_1_sqmuxa), .Q(scandata[11]));
    NOR2B state_1ms_data_1_sqmuxa_0_a2_0_0 (.A(xa_c[3]), .B(xa_c[4]), 
        .Y(state_1ms_data_1_sqmuxa_0_a2_0_net_1));
    NOR2 state_1ms_load_3_i_o2_0 (.A(N_136), .B(N_132), .Y(N_148));
    DFN1E1 \halfdata[7]  (.D(un1_GPMI_0_1[7]), .CLK(GLA), .E(
        halfdata_1_sqmuxa), .Q(halfdata[7]));
    DFN1E1 \s_acqnum[10]  (.D(un1_GPMI_0_1[10]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[10]));
    OR2 bri_datain_1_sqmuxa_0_a2_0_a2_0 (.A(N_446), .B(N_278), .Y(
        N_458));
    DFN1E1 \state_1ms_data[6]  (.D(un1_GPMI_0_1[6]), .CLK(GLA), .E(
        state_1ms_data_1_sqmuxa), .Q(state_1ms_data[6]));
    AO1A pluse_scale_RNO (.A(N_1558), .B(pluse_scale_3_0_a2_0_4), .C(
        N_215), .Y(pluse_scale_3));
    DFN1E1 \sd_sacq_data[11]  (.D(un1_GPMI_0_1[11]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[11]));
    VCC VCC_i (.Y(VCC));
    NOR2 sd_sacq_data_1_sqmuxa_0_a2_0_a2 (.A(N_451), .B(N_448), .Y(
        sd_sacq_data_1_sqmuxa));
    OA1 n_s_ctrl_RNI1LBO2 (.A(N_129), .B(n_s_ctrl_3_0_o2_0), .C(
        top_code_0_n_s_ctrl), .Y(N_217));
    MX2 \relayclose_on_RNO_0[5]  (.A(relayclose_on_c[5]), .B(
        un1_GPMI_0_1[5]), .S(relayclose_on_1_sqmuxa), .Y(N_801));
    DFN1E1 pd_pluse_load (.D(N_179), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pd_pluse_load));
    DFN1E1 \dds_configdata[15]  (.D(un1_GPMI_0_1[15]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[15]));
    NOR2A un1_xa_10_0_a2_0_a2_1 (.A(xa_c[3]), .B(N_264), .Y(
        un1_xa_10_0_a2_0_a2_1_net_1));
    NOR3B scale_rst_RNO_2 (.A(un1_state_1ms_rst_n113_35_i_a2_1), .B(
        un1_state_1ms_rst_n113_35_i_a2_0), .C(N_1558), .Y(N_210));
    DFN1E1 \pd_pluse_data[3]  (.D(un1_GPMI_0_1[3]), .CLK(GLA), .E(
        pd_pluse_data_1_sqmuxa), .Q(pd_pluse_data[3]));
    DFN1E1 \sd_sacq_data[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        sd_sacq_data_1_sqmuxa), .Q(sd_sacq_data[5]));
    MX2 noise_rst_0_0_RNILNIQ2 (.A(top_code_0_noise_rst_0), .B(
        xa_c_0_0), .S(N_164), .Y(N_792));
    OA1A state_1ms_load_RNO (.A(N_159), .B(N_136), .C(N_192), .Y(
        state_1ms_load_RNO_net_1));
    DFN1E1 \noisedata[12]  (.D(un1_GPMI_0_1[12]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[12]));
    DFN1E1 \dds_configdata[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[4]));
    DFN1E1 \sigtimedata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        sigtimedata_1_sqmuxa), .Q(sigtimedata[8]));
    NOR2B \relayclose_on_RNO[7]  (.A(N_803), .B(net_27), .Y(N_52));
    AO1C cal_load_RNO (.A(N_286), .B(cal_load_3_i_i_a2_0_0), .C(N_379), 
        .Y(N_106));
    DFN1E1 \dds_configdata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        dds_configdata_1_sqmuxa), .Q(dds_configdata[8]));
    OR3A sigrst_RNO_2 (.A(xa_c_0_7), .B(N_277), .C(xa_c_0_0), .Y(
        sigrst_3_i_a2_0_0));
    OR2 un1_state_1ms_rst_n113_43_i_a2_5 (.A(xa_c[7]), .B(xa_c[4]), .Y(
        N_232));
    DFN1 \relayclose_on[13]  (.D(N_69), .CLK(GLA), .Q(
        relayclose_on_c[13]));
    NOR3A pluseload_RNO_0 (.A(N_144_i_0), .B(N_134), .C(N_140), .Y(
        N_1565));
    DFN1E1 RAM_Rd_rst (.D(N_1544), .CLK(GLA), .E(net_27), .Q(
        top_code_0_RAM_Rd_rst));
    NOR2B \relayclose_on_RNO[0]  (.A(N_796), .B(net_27), .Y(N_95));
    DFN1E1 \s_addchoice[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        s_addchoice_1_sqmuxa), .Q(s_addchoice[2]));
    DFN1E1 \s_acqnum[2]  (.D(un1_GPMI_0_1[2]), .CLK(GLA), .E(
        s_acqnum_1_sqmuxa), .Q(s_acqnum_0[2]));
    OR3B n_rd_en_3_0_i_o2_0 (.A(N_268), .B(N_269), .C(N_229), .Y(N_290)
        );
    DFN1E1 \noisedata[8]  (.D(un1_GPMI_0_1[8]), .CLK(GLA), .E(
        noisedata_1_sqmuxa), .Q(noisedata[8]));
    DFN1E1 \scaledatain[4]  (.D(un1_GPMI_0_1[4]), .CLK(GLA), .E(
        scaledatain_1_sqmuxa), .Q(scaledatain[4]));
    AO1 scan_start_RNO_2 (.A(un1_state_1ms_rst_n113_43_i_a2_0), .B(
        un1_state_1ms_rst_n113_42_i_a2_1), .C(N_123), .Y(
        un1_state_1ms_rst_n113_42_i_0));
    DFN1 state_1ms_start (.D(N_93), .CLK(GLA), .Q(
        top_code_0_state_1ms_start));
    DFN1E1 \scaleddsdiv[5]  (.D(un1_GPMI_0_1[5]), .CLK(GLA), .E(
        scaleddsdiv_1_sqmuxa), .Q(scaleddsdiv[5]));
    MX2B pluse_lc_RNO (.A(top_code_0_pluse_lc), .B(xa_c[0]), .S(N_311), 
        .Y(N_70));
    OR3A scanchoice_RNO_0 (.A(xa_c[4]), .B(N_128), .C(N_151), .Y(N_178)
        );
    DFN1 \relayclose_on[0]  (.D(N_95), .CLK(GLA), .Q(
        relayclose_on_c[0]));
    DFN1E1 pluse_scale (.D(pluse_scale_3), .CLK(GLA), .E(net_27), .Q(
        top_code_0_pluse_scale));
    DFN1E1 sd_sacq_load (.D(N_201), .CLK(GLA), .E(net_27), .Q(
        top_code_0_sd_sacq_load));
    NOR2A cal_load_RNO_0 (.A(xa_c_0_0), .B(N_277), .Y(
        cal_load_3_i_i_a2_0_0));
    DFN1 \relayclose_on[4]  (.D(\relayclose_on_RNO[4]_net_1 ), .CLK(
        GLA), .Q(relayclose_on_c[4]));
    
endmodule


module scan_scale_sw(
       change,
       un1_top_code_0_3_0,
       ddsclkout_c,
       net_27,
       scan_scale_sw_0_s_start,
       sd_acq_en_c,
       scanstate_0_s_acq
    );
input  [1:1] change;
input  [0:0] un1_top_code_0_3_0;
input  ddsclkout_c;
input  net_27;
output scan_scale_sw_0_s_start;
input  sd_acq_en_c;
input  scanstate_0_s_acq;

    wire s_start_5, N_26, s_start_RNO_net_1, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    MX2 s_start_RNO_1 (.A(scanstate_0_s_acq), .B(sd_acq_en_c), .S(
        un1_top_code_0_3_0[0]), .Y(s_start_5));
    MX2 s_start_RNO_0 (.A(s_start_5), .B(scan_scale_sw_0_s_start), .S(
        change[1]), .Y(N_26));
    NOR2B s_start_RNO (.A(net_27), .B(N_26), .Y(s_start_RNO_net_1));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    DFN1 s_start (.D(s_start_RNO_net_1), .CLK(ddsclkout_c), .Q(
        scan_scale_sw_0_s_start));
    GND GND_i (.Y(GND));
    
endmodule


module dds_timer(
       count_2,
       count_0,
       GLA,
       dds_change_0_dds_rst,
       dds_change_0_dds_conf,
       dds_state_0_state_over
    );
output [4:0] count_2;
output [7:5] count_0;
input  GLA;
input  dds_change_0_dds_rst;
input  dds_change_0_dds_conf;
input  dds_state_0_state_over;

    wire count_0_sqmuxa_0_net_1, count_0_sqmuxa_net_1, N_17, N_23, 
        N_15, N_22, N_13, N_21, N_11, N_42, N_9, N_19, N_7, N_18, N_5, 
        count_n0, GND, VCC, GND_0, VCC_0;
    
    XA1B \count_RNO[6]  (.A(N_22), .B(count_0[6]), .C(
        count_0_sqmuxa_net_1), .Y(N_15));
    DFN1 \count[5]  (.D(N_13), .CLK(GLA), .Q(count_0[5]));
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_2[0]), .B(count_2[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_2[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_2[0]));
    XA1B \count_RNO[3]  (.A(N_19), .B(count_2[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    XA1B \count_RNO[5]  (.A(N_21), .B(count_0[5]), .C(
        count_0_sqmuxa_net_1), .Y(N_13));
    OR2B \count_RNIJ34D[0]  (.A(count_2[1]), .B(count_2[0]), .Y(N_18));
    NOR2B count_0_sqmuxa_0 (.A(dds_state_0_state_over), .B(
        dds_change_0_dds_conf), .Y(count_0_sqmuxa_0_net_1));
    NOR2B \count_RNO_0[7]  (.A(count_0[6]), .B(N_22), .Y(N_23));
    XA1B \count_RNO[7]  (.A(N_23), .B(count_0[7]), .C(
        count_0_sqmuxa_net_1), .Y(N_17));
    NOR2A \count_RNIEBMJ[2]  (.A(count_2[2]), .B(N_18), .Y(N_19));
    GND GND_i (.Y(GND));
    AOI1 \count_RNO_0[4]  (.A(count_2[3]), .B(N_19), .C(count_2[4]), 
        .Y(N_42));
    NOR2B \count_RNI5RD71[5]  (.A(count_0[5]), .B(N_21), .Y(N_22));
    XA1C \count_RNO[2]  (.A(N_18), .B(count_2[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR2B count_0_sqmuxa (.A(count_0_sqmuxa_0_net_1), .B(
        dds_change_0_dds_rst), .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR3 \count_RNO[4]  (.A(N_42), .B(count_0_sqmuxa_net_1), .C(N_21), 
        .Y(N_11));
    NOR3C \count_RNI77R01[4]  (.A(N_19), .B(count_2[3]), .C(count_2[4])
        , .Y(N_21));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_2[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_2[4]));
    NOR2 \count_RNO[0]  (.A(count_2[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[6]  (.D(N_15), .CLK(GLA), .Q(count_0[6]));
    DFN1 \count[7]  (.D(N_17), .CLK(GLA), .Q(count_0[7]));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_2[2]));
    
endmodule


module dds_state(
       i_2,
       dds_configdata,
       i_RNIV2B7,
       ddsreset_c,
       ddsdata_c,
       ddsfqud_c,
       ddswclk_c,
       GLA,
       dds_change_0_dds_rst,
       dds_state_0_state_over,
       top_code_0_dds_choice,
       top_code_0_dds_load
    );
input  [3:1] i_2;
input  [15:0] dds_configdata;
input  [0:0] i_RNIV2B7;
output ddsreset_c;
output ddsdata_c;
output ddsfqud_c;
output ddswclk_c;
input  GLA;
input  dds_change_0_dds_rst;
output dds_state_0_state_over;
input  top_code_0_dds_choice;
input  top_code_0_dds_load;

    wire N_540_1, N_540_0, N_572_1, N_572_0, para_1_sqmuxa_1_0, 
        w_clk_reg_net_1, \para_9_i_0[7] , N_436, \para_9_i_0[15] , 
        N_440, \para_9_i_0[20] , N_444, \para_9_i_0[21] , N_448, 
        \para_9_i_0[22] , N_452, \para_9_i_0[30] , N_456, 
        \para_9_i_0[1] , N_474, \para_9_i_0[2] , N_478, 
        \para_9_i_0[3] , N_482, \para_9_i_0[4] , N_486, 
        \para_9_i_0[17] , N_343, \para_9_i_0[18] , N_347, 
        \para_9_i_0[19] , N_351, \para_9_i_0[31] , N_355, 
        \para_9_i_0[12] , N_365, \para_9_i_0[13] , N_369, 
        \para_9_i_0[14] , N_373, \para_9_i_0[27] , N_380, 
        \para_9_i_0[28] , N_387, \para_9_i_0[29] , N_391, 
        \para_9_i_0[5] , N_405, \para_9_i_0[6] , N_489, 
        \para_9_i_0[8] , N_493, \para_9_i_0[9] , N_497, 
        \para_9_i_0[10] , N_501, \para_9_i_0[11] , N_505, 
        \para_9_i_0[16] , N_509, \para_9_i_0[23] , N_513, 
        \para_9_i_0[24] , N_517, \para_9_i_0[25] , N_521, 
        \para_9_i_0[26] , N_525, \para_9_i_0[32] , N_529, N_167, N_528, 
        N_527, N_165, N_524, N_523, N_163, N_520, N_519, N_161, N_516, 
        N_515, N_159, N_512, N_511, N_157, N_508, N_507, N_155, N_504, 
        N_503, N_153, N_500, N_499, N_151, N_496, N_495, N_149, N_492, 
        N_491, N_147, N_488, N_487, N_145, N_396, N_394, N_143, N_390, 
        N_389, N_141, N_386, N_384, N_139, N_378, N_376, N_137, N_372, 
        N_371, N_135, N_368, N_367, N_133, N_364, N_363, N_128, N_354, 
        N_353, N_126, N_350, N_349, N_124, N_346, N_345, N_122, N_342, 
        N_341, N_120, N_485, N_484, N_46, N_481, N_480, N_44, N_477, 
        N_476, N_42, N_473, N_472, N_15, N_455, N_454, N_13, N_451, 
        N_450, N_11, N_447, N_446, N_9, N_443, N_442, N_7, N_439, 
        N_438, N_5, N_435, N_434, N_37, N_466, \para[0]_net_1 , N_238, 
        N_539, \cs[8]_net_1 , \cs[7]_net_1 , para_1_sqmuxa_1, 
        \para[7]_net_1 , \para[8]_net_1 , \para_reg[7]_net_1 , 
        \para[15]_net_1 , \para[16]_net_1 , \para_reg[15]_net_1 , 
        \para[20]_net_1 , \para[21]_net_1 , \para_reg[20]_net_1 , 
        \para[22]_net_1 , \para_reg[21]_net_1 , \para[23]_net_1 , 
        \para_reg[22]_net_1 , \para[30]_net_1 , \para[31]_net_1 , 
        \para_reg[30]_net_1 , \cs_RNO_1[3] , N_242, \cs_RNO_0[4] , 
        \cs[3]_net_1 , \cs_RNO_0[6] , \cs[5]_net_1 , \cs_RNO_0[7] , 
        N_241, \cs_RNO[8]_net_1 , w_clk_RNO_net_1, fq_ud_RNO_net_1, 
        fq_ud_reg_net_1, N_239, \cs[4]_net_1 , reset_RNO_net_1, 
        \cs[1]_net_1 , N_470, \para[1]_net_1 , \para[2]_net_1 , 
        \para_reg[1]_net_1 , \para[3]_net_1 , \para_reg[2]_net_1 , 
        \para[4]_net_1 , \para_reg[3]_net_1 , \para[5]_net_1 , 
        \para_reg[4]_net_1 , \para[17]_net_1 , \para[18]_net_1 , 
        \para_reg[17]_net_1 , \para[19]_net_1 , \para_reg[18]_net_1 , 
        \para_reg[19]_net_1 , \para[32]_net_1 , \para_reg[31]_net_1 , 
        N_357, \para[34]_net_1 , N_359, \para[35]_net_1 , N_361, 
        \para[36]_net_1 , \para[12]_net_1 , \para[13]_net_1 , 
        \para_reg[12]_net_1 , \para[14]_net_1 , \para_reg[13]_net_1 , 
        \para_reg[14]_net_1 , \para[27]_net_1 , \para[28]_net_1 , 
        \para_reg[27]_net_1 , \para[29]_net_1 , \para_reg[28]_net_1 , 
        \para_reg[29]_net_1 , \para[6]_net_1 , \para_reg[5]_net_1 , 
        \para_reg[6]_net_1 , \para[9]_net_1 , \para_reg[8]_net_1 , 
        \para[10]_net_1 , \para_reg[9]_net_1 , \para[11]_net_1 , 
        \para_reg[10]_net_1 , \para_reg[11]_net_1 , 
        \para_reg[16]_net_1 , \para[24]_net_1 , \para_reg[23]_net_1 , 
        \para[25]_net_1 , \para_reg[24]_net_1 , \para[26]_net_1 , 
        \para_reg[25]_net_1 , \para_reg[26]_net_1 , \para[33]_net_1 , 
        \para_reg[32]_net_1 , \para_9[36] , N_19, N_243, N_240, 
        \cs_RNO_0[5] , fq_ud_reg_RNO_net_1, w_clk_reg_RNO_net_1, 
        \cs_RNO_0[1]_net_1 , \cs_i[0]_net_1 , N_244, 
        state_over_RNO_net_1, \para_9[0] , \para_9[33] , \para_9[34] , 
        \para_9[35] , \cs[6]_net_1 , \cs[2]_net_1 , N_572, N_540, GND, 
        VCC, GND_0, VCC_0;
    
    NOR2 \para_RNO_1[8]  (.A(\para[8]_net_1 ), .B(N_572_1), .Y(N_491));
    NOR3A \para_RNO_0[29]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[30]_net_1 ), .Y(N_390));
    NOR3 \para_RNO[7]  (.A(N_435), .B(N_434), .C(\para_9_i_0[7] ), .Y(
        N_5));
    NOR3 \para_RNO[5]  (.A(N_396), .B(N_394), .C(\para_9_i_0[5] ), .Y(
        N_145));
    DFN1E0 \para_reg[2]  (.D(dds_configdata[1]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[2]_net_1 ));
    NOR2 \para_RNO_1[10]  (.A(\para[10]_net_1 ), .B(N_572_1), .Y(N_499)
        );
    NOR3 \para_RNO[20]  (.A(N_443), .B(N_442), .C(\para_9_i_0[20] ), 
        .Y(N_9));
    DFN1E0 \para[35]  (.D(\para_9[35] ), .CLK(GLA), .E(para_1_sqmuxa_1)
        , .Q(\para[35]_net_1 ));
    DFN1E0 \para[21]  (.D(N_11), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[21]_net_1 ));
    NOR3A \para_RNO_0[6]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[7]_net_1 ), .Y(N_488));
    NOR3A \para_RNO_0[26]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[27]_net_1 ), .Y(N_524));
    OR2A para_reg_18_e_0 (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_540_0));
    AO1D \para_RNO_2[22]  (.A(dds_configdata[5]), .B(N_572_0), .C(
        N_452), .Y(\para_9_i_0[22] ));
    NOR3 \para_RNO[16]  (.A(N_508), .B(N_507), .C(\para_9_i_0[16] ), 
        .Y(N_157));
    DFN1 state_over (.D(state_over_RNO_net_1), .CLK(GLA), .Q(
        dds_state_0_state_over));
    NOR2B \cs_RNO[4]  (.A(\cs[3]_net_1 ), .B(N_238), .Y(\cs_RNO_0[4] ));
    DFN1E0 \para[22]  (.D(N_13), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[22]_net_1 ));
    NOR2 \para_RNO_1[18]  (.A(\para[18]_net_1 ), .B(N_540_1), .Y(N_345)
        );
    NOR3A \para_RNO_0[23]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[24]_net_1 ), .Y(N_512));
    DFN1E0 \para[30]  (.D(N_15), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[30]_net_1 ));
    NOR3A \para_RNO_0[8]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[9]_net_1 ), .Y(N_492));
    NOR3A \para_RNO_0[25]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[26]_net_1 ), .Y(N_520));
    AO1D \para_RNO_2[2]  (.A(dds_configdata[1]), .B(N_540_0), .C(N_478)
        , .Y(\para_9_i_0[2] ));
    OR3B \para_RNO_0[33]  (.A(i_RNIV2B7[0]), .B(\para[34]_net_1 ), .C(
        top_code_0_dds_load), .Y(N_357));
    AO1D \para_RNO_2[29]  (.A(dds_configdata[12]), .B(N_572_0), .C(
        N_391), .Y(\para_9_i_0[29] ));
    OR3B \para_RNO_0[35]  (.A(i_RNIV2B7[0]), .B(\para[36]_net_1 ), .C(
        top_code_0_dds_load), .Y(N_361));
    DFN1 \cs[4]  (.D(\cs_RNO_0[4] ), .CLK(GLA), .Q(\cs[4]_net_1 ));
    NOR2B \cs_RNICV1B[6]  (.A(i_2[3]), .B(\cs[6]_net_1 ), .Y(N_241));
    NOR3 \para_RNO[6]  (.A(N_488), .B(N_487), .C(\para_9_i_0[6] ), .Y(
        N_147));
    NOR3 \para_RNO_3[11]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[11]_net_1 ), .Y(N_505));
    NOR3A \para_RNO_0[11]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[12]_net_1 ), .Y(N_504));
    AO1D \para_RNO_2[31]  (.A(dds_configdata[14]), .B(N_572_0), .C(
        N_355), .Y(\para_9_i_0[31] ));
    DFN1E0 \para[19]  (.D(N_126), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[19]_net_1 ));
    NOR3 \para_RNO_3[22]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[22]_net_1 ), .Y(N_452));
    NOR2 \para_RNO_1[32]  (.A(\para[32]_net_1 ), .B(N_540_1), .Y(N_527)
        );
    AO1D \para_RNO_2[11]  (.A(dds_configdata[10]), .B(N_540_0), .C(
        N_505), .Y(\para_9_i_0[11] ));
    OR2A \cs_RNO_1[2]  (.A(\cs[2]_net_1 ), .B(i_2[2]), .Y(N_240));
    NOR2B cs4_i_i_o2 (.A(dds_change_0_dds_rst), .B(i_RNIV2B7[0]), .Y(
        N_238));
    DFN1E0 \para_reg[6]  (.D(dds_configdata[5]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[6]_net_1 ));
    NOR3 \para_RNO_3[17]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[17]_net_1 ), .Y(N_343));
    NOR3A \para_RNO_0[17]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[18]_net_1 ), .Y(N_342));
    AO1D \para_RNO_2[9]  (.A(dds_configdata[8]), .B(N_540_0), .C(N_497)
        , .Y(\para_9_i_0[9] ));
    AO1D \para_RNO_2[26]  (.A(dds_configdata[9]), .B(N_572_0), .C(
        N_525), .Y(\para_9_i_0[26] ));
    NOR2 \para_RNO_1[21]  (.A(\para[21]_net_1 ), .B(N_540_0), .Y(N_446)
        );
    AO1D \para_RNO_2[17]  (.A(dds_configdata[0]), .B(N_572_0), .C(
        N_343), .Y(\para_9_i_0[17] ));
    DFN1E0 \para[27]  (.D(N_139), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[27]_net_1 ));
    NOR3 \para_RNO_3[14]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[14]_net_1 ), .Y(N_373));
    NOR3A \para_RNO_0[14]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[15]_net_1 ), .Y(N_372));
    NOR2B \cs_RNI7R1B[2]  (.A(i_2[2]), .B(\cs[2]_net_1 ), .Y(N_242));
    DFN1E0 \para[23]  (.D(N_159), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[23]_net_1 ));
    NOR2 \para_RNO_1[27]  (.A(\para[27]_net_1 ), .B(N_540_1), .Y(N_376)
        );
    NOR3 \para_RNO_3[29]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[29]_net_1 ), .Y(N_391));
    AO1D \para_RNO_2[14]  (.A(dds_configdata[13]), .B(N_540_0), .C(
        N_373), .Y(\para_9_i_0[14] ));
    DFN1 \cs[3]  (.D(\cs_RNO_1[3] ), .CLK(GLA), .Q(\cs[3]_net_1 ));
    AO1D \para_RNO_2[23]  (.A(dds_configdata[6]), .B(N_572_0), .C(
        N_513), .Y(\para_9_i_0[23] ));
    NOR2 \para_RNO_1[24]  (.A(\para[24]_net_1 ), .B(N_540_1), .Y(N_515)
        );
    AO1D \para_RNO_2[25]  (.A(dds_configdata[8]), .B(N_572_0), .C(
        N_521), .Y(\para_9_i_0[25] ));
    AO1C \para_RNO[33]  (.A(N_540_1), .B(\para[33]_net_1 ), .C(N_357), 
        .Y(\para_9[33] ));
    OA1 fq_ud_reg_RNO (.A(N_241), .B(\cs[3]_net_1 ), .C(N_238), .Y(
        fq_ud_reg_RNO_net_1));
    NOR2B w_clk_RNO (.A(w_clk_reg_net_1), .B(N_238), .Y(
        w_clk_RNO_net_1));
    OA1 \cs_RNO[5]  (.A(N_239), .B(\cs[4]_net_1 ), .C(N_238), .Y(
        \cs_RNO_0[5] ));
    NOR3 \para_RNO_3[4]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[4]_net_1 ), .Y(N_486));
    NOR3 \para_RNO[14]  (.A(N_372), .B(N_371), .C(\para_9_i_0[14] ), 
        .Y(N_137));
    NOR3 \para_RNO_3[32]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[32]_net_1 ), .Y(N_529));
    NOR3A \para_RNO_0[4]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[5]_net_1 ), .Y(N_485));
    NOR3 \para_RNO_3[26]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[26]_net_1 ), .Y(N_525));
    NOR3 \para_RNO[11]  (.A(N_504), .B(N_503), .C(\para_9_i_0[11] ), 
        .Y(N_155));
    NOR3 \para_RNO[22]  (.A(N_451), .B(N_450), .C(\para_9_i_0[22] ), 
        .Y(N_13));
    NOR3 \para_RNO_3[10]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[10]_net_1 ), .Y(N_501));
    NOR3A \para_RNO_0[10]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[11]_net_1 ), .Y(N_500));
    OR2A \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_2[1]), .Y(N_244));
    AO1D \para_RNO_2[30]  (.A(dds_configdata[13]), .B(N_572_0), .C(
        N_456), .Y(\para_9_i_0[30] ));
    DFN1E0 \para[11]  (.D(N_155), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[11]_net_1 ));
    AO1D \para_RNO_2[10]  (.A(dds_configdata[9]), .B(N_540_0), .C(
        N_501), .Y(\para_9_i_0[10] ));
    DFN1 \cs[1]  (.D(\cs_RNO_0[1]_net_1 ), .CLK(GLA), .Q(\cs[1]_net_1 )
        );
    DFN1E0 \para[26]  (.D(N_165), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[26]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1 data (.D(N_37), .CLK(GLA), .Q(ddsdata_c));
    AO1D \para_RNO_2[6]  (.A(dds_configdata[5]), .B(N_540_0), .C(N_489)
        , .Y(\para_9_i_0[6] ));
    NOR2 \para_RNO_1[20]  (.A(\para[20]_net_1 ), .B(N_540_0), .Y(N_442)
        );
    NOR3A \para_RNO_0[21]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[22]_net_1 ), .Y(N_447));
    NOR3 \para_RNO_3[23]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[23]_net_1 ), .Y(N_513));
    NOR3A \para_RNO_0[31]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[32]_net_1 ), .Y(N_354));
    DFN1 reset (.D(reset_RNO_net_1), .CLK(GLA), .Q(ddsreset_c));
    NOR3 \para_RNO_3[25]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[25]_net_1 ), .Y(N_521));
    DFN1E0 \para[12]  (.D(N_133), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[12]_net_1 ));
    DFN1 \cs_i[0]  (.D(N_238), .CLK(GLA), .Q(\cs_i[0]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR3A \para_RNO_0[27]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[28]_net_1 ), .Y(N_378));
    NOR3A \para_RNO_0[7]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[8]_net_1 ), .Y(N_435));
    NOR3 \para_RNO_3[18]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[18]_net_1 ), .Y(N_347));
    NOR3A \para_RNO_0[18]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[19]_net_1 ), .Y(N_346));
    DFN1E0 \para_reg[3]  (.D(dds_configdata[2]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[3]_net_1 ));
    DFN1 w_clk (.D(w_clk_RNO_net_1), .CLK(GLA), .Q(ddswclk_c));
    NOR2B \cs_RNO[7]  (.A(N_241), .B(N_238), .Y(\cs_RNO_0[7] ));
    NOR3A \para_RNO_0[24]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[25]_net_1 ), .Y(N_516));
    AO1D \para_RNO_2[18]  (.A(dds_configdata[1]), .B(N_572_0), .C(
        N_347), .Y(\para_9_i_0[18] ));
    NOR3 \para_RNO[25]  (.A(N_520), .B(N_519), .C(\para_9_i_0[25] ), 
        .Y(N_163));
    NOR3 \para_RNO_3[6]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[6]_net_1 ), .Y(N_489));
    OR3B \para_RNO_0[34]  (.A(i_RNIV2B7[0]), .B(\para[35]_net_1 ), .C(
        top_code_0_dds_load), .Y(N_359));
    NOR2 \para_RNO_1[28]  (.A(\para[28]_net_1 ), .B(N_540_1), .Y(N_384)
        );
    DFN1E0 \para_reg[27]  (.D(dds_configdata[10]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[27]_net_1 ));
    DFN1E0 \para_reg[29]  (.D(dds_configdata[12]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[29]_net_1 ));
    DFN1E0 \para[3]  (.D(N_46), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[3]_net_1 ));
    NOR3 \para_RNO_3[7]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[7]_net_1 ), .Y(N_436));
    DFN1E0 \para[5]  (.D(N_145), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[5]_net_1 ));
    NOR2B \cs_RNO[3]  (.A(N_242), .B(N_238), .Y(\cs_RNO_1[3] ));
    AO1D \para_RNO_2[21]  (.A(dds_configdata[4]), .B(N_572_0), .C(
        N_448), .Y(\para_9_i_0[21] ));
    DFN1E0 \para_reg[17]  (.D(dds_configdata[0]), .CLK(GLA), .E(
        N_572_1), .Q(\para_reg[17]_net_1 ));
    DFN1E0 \para[17]  (.D(N_122), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[17]_net_1 ));
    DFN1E0 \para_reg[19]  (.D(dds_configdata[2]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[19]_net_1 ));
    NOR3A \para_RNO_0[20]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[21]_net_1 ), .Y(N_443));
    AO1C \para_RNO[0]  (.A(N_572_1), .B(\para[0]_net_1 ), .C(N_470), 
        .Y(\para_9[0] ));
    NOR3A \para_RNO_0[2]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[3]_net_1 ), .Y(N_477));
    DFN1E0 \para[13]  (.D(N_135), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[13]_net_1 ));
    NOR3A \para_RNO_0[30]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[31]_net_1 ), .Y(N_455));
    NOR3 \para_RNO[26]  (.A(N_524), .B(N_523), .C(\para_9_i_0[26] ), 
        .Y(N_165));
    AOI1B \cs_RNO[1]  (.A(\cs_i[0]_net_1 ), .B(N_244), .C(N_238), .Y(
        \cs_RNO_0[1]_net_1 ));
    AO1D \para_RNO_2[27]  (.A(dds_configdata[10]), .B(N_572_0), .C(
        N_380), .Y(\para_9_i_0[27] ));
    VCC VCC_i (.Y(VCC));
    DFN1E0 \para_reg[8]  (.D(dds_configdata[7]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[8]_net_1 ));
    DFN1E0 \para_reg[24]  (.D(dds_configdata[7]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[24]_net_1 ));
    AO1D \para_RNO_2[24]  (.A(dds_configdata[7]), .B(N_572_0), .C(
        N_517), .Y(\para_9_i_0[24] ));
    DFN1E0 \para[28]  (.D(N_141), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[28]_net_1 ));
    OR2B \cs_RNO_0[2]  (.A(i_2[1]), .B(\cs[1]_net_1 ), .Y(N_243));
    DFN1E0 \para[9]  (.D(N_151), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[9]_net_1 ));
    NOR3A \para_RNO_0[5]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[6]_net_1 ), .Y(N_396));
    NOR3A \para_RNO_0[28]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[29]_net_1 ), .Y(N_386));
    NOR3 \para_RNO[18]  (.A(N_346), .B(N_345), .C(\para_9_i_0[18] ), 
        .Y(N_124));
    DFN1E0 \para_reg[5]  (.D(dds_configdata[4]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[5]_net_1 ));
    DFN1E0 \para_reg[25]  (.D(dds_configdata[8]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[25]_net_1 ));
    NOR3 \para_RNO_3[21]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[21]_net_1 ), .Y(N_448));
    DFN1E0 \para_reg[14]  (.D(dds_configdata[13]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[14]_net_1 ));
    DFN1E0 \para[31]  (.D(N_128), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[31]_net_1 ));
    NOR3 \para_RNO_3[2]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[2]_net_1 ), .Y(N_478));
    NOR2 \para_RNO_1[31]  (.A(\para[31]_net_1 ), .B(N_540_1), .Y(N_353)
        );
    NOR3 \para_RNO[30]  (.A(N_455), .B(N_454), .C(\para_9_i_0[30] ), 
        .Y(N_15));
    DFN1E0 \para[16]  (.D(N_157), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[16]_net_1 ));
    NOR3 \para_RNO_3[27]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[27]_net_1 ), .Y(N_380));
    AO1D \para_RNO_2[20]  (.A(dds_configdata[3]), .B(N_572_0), .C(
        N_444), .Y(\para_9_i_0[20] ));
    DFN1E0 \para_reg[15]  (.D(dds_configdata[14]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[15]_net_1 ));
    DFN1E0 \para[32]  (.D(N_167), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[32]_net_1 ));
    NOR3 \para_RNO_3[24]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[24]_net_1 ), .Y(N_517));
    NOR3 \para_RNO_3[3]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[3]_net_1 ), .Y(N_482));
    DFN1E0 \para[4]  (.D(N_120), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[4]_net_1 ));
    NOR3 \para_RNO[19]  (.A(N_350), .B(N_349), .C(\para_9_i_0[19] ), 
        .Y(N_126));
    OR2B para_reg_34_e_1 (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_572_1));
    DFN1 fq_ud_reg (.D(fq_ud_reg_RNO_net_1), .CLK(GLA), .Q(
        fq_ud_reg_net_1));
    NOR3 \para_RNO_3[31]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[31]_net_1 ), .Y(N_355));
    AO1D \para_RNO_2[28]  (.A(dds_configdata[11]), .B(N_572_0), .C(
        N_387), .Y(\para_9_i_0[28] ));
    NOR3 \para_RNO[13]  (.A(N_368), .B(N_367), .C(\para_9_i_0[13] ), 
        .Y(N_135));
    DFN1E0 \para[24]  (.D(N_161), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[24]_net_1 ));
    NOR3 \para_RNO[24]  (.A(N_516), .B(N_515), .C(\para_9_i_0[24] ), 
        .Y(N_161));
    NOR3 \para_RNO_3[20]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[20]_net_1 ), .Y(N_444));
    NOR3 \para_RNO[21]  (.A(N_447), .B(N_446), .C(\para_9_i_0[21] ), 
        .Y(N_11));
    NOR2B fq_ud_RNO (.A(fq_ud_reg_net_1), .B(N_238), .Y(
        fq_ud_RNO_net_1));
    NOR2 \para_RNO_1[30]  (.A(\para[30]_net_1 ), .B(N_540_1), .Y(N_454)
        );
    OR3B \para_RNO_0[0]  (.A(i_RNIV2B7[0]), .B(\para[1]_net_1 ), .C(
        top_code_0_dds_load), .Y(N_470));
    NOR3 \para_RNO_3[5]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[5]_net_1 ), .Y(N_405));
    DFN1E0 \para[33]  (.D(\para_9[33] ), .CLK(GLA), .E(para_1_sqmuxa_1)
        , .Q(\para[33]_net_1 ));
    NOR3 \para_RNO[3]  (.A(N_481), .B(N_480), .C(\para_9_i_0[3] ), .Y(
        N_46));
    NOR3 \para_RNO_3[1]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[1]_net_1 ), .Y(N_474));
    AO1D \para_RNO_2[8]  (.A(dds_configdata[7]), .B(N_540_0), .C(N_493)
        , .Y(\para_9_i_0[8] ));
    NOR3 \para_RNO_3[28]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[28]_net_1 ), .Y(N_387));
    DFN1 \cs[7]  (.D(\cs_RNO_0[7] ), .CLK(GLA), .Q(\cs[7]_net_1 ));
    DFN1E0 \para[18]  (.D(N_124), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[18]_net_1 ));
    OR2B para_reg_34_e (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_572));
    AO1D \para_RNO_2[7]  (.A(dds_configdata[6]), .B(N_540_0), .C(N_436)
        , .Y(\para_9_i_0[7] ));
    DFN1 \cs[6]  (.D(\cs_RNO_0[6] ), .CLK(GLA), .Q(\cs[6]_net_1 ));
    NOR3 \para_RNO_3[30]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[30]_net_1 ), .Y(N_456));
    NOR3 \para_RNO[17]  (.A(N_342), .B(N_341), .C(\para_9_i_0[17] ), 
        .Y(N_122));
    NOR3 \para_RNO[32]  (.A(N_528), .B(N_527), .C(\para_9_i_0[32] ), 
        .Y(N_167));
    NOR2 \para_RNO_1[9]  (.A(\para[9]_net_1 ), .B(N_572_1), .Y(N_495));
    DFN1E0 \para[1]  (.D(N_42), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[1]_net_1 ));
    DFN1E0 \para[36]  (.D(\para_9[36] ), .CLK(GLA), .E(para_1_sqmuxa_1)
        , .Q(\para[36]_net_1 ));
    DFN1E0 \para[6]  (.D(N_147), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[6]_net_1 ));
    NOR2 \para_RNO_1[12]  (.A(\para[12]_net_1 ), .B(N_572_1), .Y(N_363)
        );
    OR2A para_reg_18_e_1 (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_540_1));
    NOR3A \para_RNO_0[9]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[10]_net_1 ), .Y(N_496));
    DFN1E0 \para[25]  (.D(N_163), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[25]_net_1 ));
    AOI1B \cs_RNO[2]  (.A(N_243), .B(N_240), .C(N_238), .Y(N_19));
    GND GND_i_0 (.Y(GND_0));
    AO1D \para_RNO_2[4]  (.A(dds_configdata[3]), .B(N_540_0), .C(N_486)
        , .Y(\para_9_i_0[4] ));
    DFN1E0 \para_reg[31]  (.D(dds_configdata[14]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[31]_net_1 ));
    DFN1E0 \para_reg[30]  (.D(dds_configdata[13]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[30]_net_1 ));
    DFN1E0 \para_reg[28]  (.D(dds_configdata[11]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[28]_net_1 ));
    NOR3 \para_RNO[2]  (.A(N_477), .B(N_476), .C(\para_9_i_0[2] ), .Y(
        N_44));
    DFN1 w_clk_reg (.D(w_clk_reg_RNO_net_1), .CLK(GLA), .Q(
        w_clk_reg_net_1));
    DFN1 \cs[8]  (.D(\cs_RNO[8]_net_1 ), .CLK(GLA), .Q(\cs[8]_net_1 ));
    DFN1E0 \para[8]  (.D(N_149), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[8]_net_1 ));
    NOR2 \para_RNO_1[3]  (.A(\para[3]_net_1 ), .B(N_572_1), .Y(N_480));
    NOR3 \para_RNO_3[9]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[9]_net_1 ), .Y(N_497));
    NOR2 \para_RNO_1[19]  (.A(\para[19]_net_1 ), .B(N_540_1), .Y(N_349)
        );
    AO1C \para_RNO[35]  (.A(N_540_1), .B(\para[35]_net_1 ), .C(N_361), 
        .Y(\para_9[35] ));
    NOR3 \para_RNO[4]  (.A(N_485), .B(N_484), .C(\para_9_i_0[4] ), .Y(
        N_120));
    NOR2 \para_RNO_1[1]  (.A(\para[1]_net_1 ), .B(N_572_1), .Y(N_472));
    DFN1E0 \para_reg[18]  (.D(dds_configdata[1]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[18]_net_1 ));
    DFN1E0 \para_reg[32]  (.D(dds_configdata[15]), .CLK(GLA), .E(N_572)
        , .Q(\para_reg[32]_net_1 ));
    DFN1E0 \para[20]  (.D(N_9), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[20]_net_1 ));
    DFN1E0 \para[14]  (.D(N_137), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[14]_net_1 ));
    NOR3 \para_RNO[28]  (.A(N_386), .B(N_384), .C(\para_9_i_0[28] ), 
        .Y(N_141));
    NOR2 \para_RNO_1[16]  (.A(\para[16]_net_1 ), .B(N_572_1), .Y(N_507)
        );
    NOR3 \para_RNO[10]  (.A(N_500), .B(N_499), .C(\para_9_i_0[10] ), 
        .Y(N_153));
    NOR2 \cs_RNIN0D7[7]  (.A(\cs[8]_net_1 ), .B(\cs[7]_net_1 ), .Y(
        N_539));
    DFN1 \cs[2]  (.D(N_19), .CLK(GLA), .Q(\cs[2]_net_1 ));
    NOR2 \para_RNO_1[2]  (.A(\para[2]_net_1 ), .B(N_572_1), .Y(N_476));
    DFN1E0 \para_reg[23]  (.D(dds_configdata[6]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[23]_net_1 ));
    NOR3A w_clk_reg_RNIC4AH_0 (.A(i_RNIV2B7[0]), .B(
        top_code_0_dds_load), .C(w_clk_reg_net_1), .Y(para_1_sqmuxa_1));
    NOR2A \para_RNO[36]  (.A(\para[36]_net_1 ), .B(N_540_1), .Y(
        \para_9[36] ));
    DFN1E0 \para[7]  (.D(N_5), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[7]_net_1 ));
    NOR2 \para_RNO_1[13]  (.A(\para[13]_net_1 ), .B(N_572_1), .Y(N_367)
        );
    NOR3A \para_RNO_0[3]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[4]_net_1 ), .Y(N_481));
    DFN1E0 \para[0]  (.D(\para_9[0] ), .CLK(GLA), .E(para_1_sqmuxa_1_0)
        , .Q(\para[0]_net_1 ));
    NOR2 \para_RNO_1[15]  (.A(\para[15]_net_1 ), .B(N_572_1), .Y(N_438)
        );
    NOR3 \para_RNO[1]  (.A(N_473), .B(N_472), .C(\para_9_i_0[1] ), .Y(
        N_42));
    DFN1E0 \para_reg[13]  (.D(dds_configdata[12]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[13]_net_1 ));
    NOR3 \para_RNO[29]  (.A(N_390), .B(N_389), .C(\para_9_i_0[29] ), 
        .Y(N_143));
    DFN1E0 \para_reg[26]  (.D(dds_configdata[9]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[26]_net_1 ));
    DFN1E0 \para_reg[4]  (.D(dds_configdata[3]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[4]_net_1 ));
    NOR3C data_RNO (.A(N_466), .B(\para[0]_net_1 ), .C(N_238), .Y(N_37)
        );
    DFN1E0 \para_reg[21]  (.D(dds_configdata[4]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[21]_net_1 ));
    DFN1E0 \para_reg[20]  (.D(dds_configdata[3]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[20]_net_1 ));
    NOR2 \para_RNO_1[5]  (.A(\para[5]_net_1 ), .B(N_572_1), .Y(N_394));
    NOR3 \para_RNO[23]  (.A(N_512), .B(N_511), .C(\para_9_i_0[23] ), 
        .Y(N_159));
    NOR2 \para_RNO_1[7]  (.A(\para[7]_net_1 ), .B(N_572_0), .Y(N_434));
    NOR3 \para_RNO_3[8]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[8]_net_1 ), .Y(N_493));
    NOR3 \para_RNO_3[12]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[12]_net_1 ), .Y(N_365));
    NOR3A \para_RNO_0[12]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[13]_net_1 ), .Y(N_364));
    DFN1E0 \para_reg[16]  (.D(dds_configdata[15]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[16]_net_1 ));
    NOR3A w_clk_reg_RNIC4AH (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(w_clk_reg_net_1), .Y(para_1_sqmuxa_1_0));
    AO1D \para_RNO_2[32]  (.A(dds_configdata[15]), .B(N_572_0), .C(
        N_529), .Y(\para_9_i_0[32] ));
    DFN1E0 \para_reg[11]  (.D(dds_configdata[10]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[11]_net_1 ));
    DFN1E0 \para_reg[10]  (.D(dds_configdata[9]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[10]_net_1 ));
    AO1D \para_RNO_2[12]  (.A(dds_configdata[11]), .B(N_540_0), .C(
        N_365), .Y(\para_9_i_0[12] ));
    DFN1E0 \para_reg[22]  (.D(dds_configdata[5]), .CLK(GLA), .E(N_572), 
        .Q(\para_reg[22]_net_1 ));
    DFN1E0 \para[15]  (.D(N_7), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[15]_net_1 ));
    NOR2B reset_RNO (.A(\cs[1]_net_1 ), .B(N_238), .Y(reset_RNO_net_1));
    NOR2 \para_RNO_1[22]  (.A(\para[22]_net_1 ), .B(N_540_1), .Y(N_450)
        );
    OA1 w_clk_reg_RNO (.A(N_242), .B(\cs[5]_net_1 ), .C(N_238), .Y(
        w_clk_reg_RNO_net_1));
    NOR2A \cs_RNO[8]  (.A(N_238), .B(N_539), .Y(\cs_RNO[8]_net_1 ));
    DFN1E0 \para_reg[7]  (.D(dds_configdata[6]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[7]_net_1 ));
    NOR3 \para_RNO_3[19]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[19]_net_1 ), .Y(N_351));
    NOR3A \para_RNO_0[19]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[20]_net_1 ), .Y(N_350));
    NOR2A \cs_RNICV1B_0[6]  (.A(\cs[6]_net_1 ), .B(i_2[3]), .Y(N_239));
    DFN1 \cs[5]  (.D(\cs_RNO_0[5] ), .CLK(GLA), .Q(\cs[5]_net_1 ));
    DFN1E0 \para_reg[1]  (.D(dds_configdata[0]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[1]_net_1 ));
    NOR2 \para_RNO_1[6]  (.A(\para[6]_net_1 ), .B(N_572_1), .Y(N_487));
    NOR3A \para_RNO_0[1]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[2]_net_1 ), .Y(N_473));
    DFN1E0 \para_reg[12]  (.D(dds_configdata[11]), .CLK(GLA), .E(N_540)
        , .Q(\para_reg[12]_net_1 ));
    AO1D \para_RNO_2[19]  (.A(dds_configdata[2]), .B(N_572_0), .C(
        N_351), .Y(\para_9_i_0[19] ));
    DFN1E0 \para[34]  (.D(\para_9[34] ), .CLK(GLA), .E(para_1_sqmuxa_1)
        , .Q(\para[34]_net_1 ));
    AO1D \para_RNO_2[3]  (.A(dds_configdata[2]), .B(N_540_0), .C(N_482)
        , .Y(\para_9_i_0[3] ));
    NOR2 \para_RNO_1[29]  (.A(\para[29]_net_1 ), .B(N_540_1), .Y(N_389)
        );
    DFN1E0 \para[10]  (.D(N_153), .CLK(GLA), .E(para_1_sqmuxa_1_0), .Q(
        \para[10]_net_1 ));
    AO1C \para_RNO[34]  (.A(N_540_1), .B(\para[34]_net_1 ), .C(N_359), 
        .Y(\para_9[34] ));
    AO1D \para_RNO_2[1]  (.A(dds_configdata[0]), .B(N_540_0), .C(N_474)
        , .Y(\para_9_i_0[1] ));
    NOR3 \para_RNO[27]  (.A(N_378), .B(N_376), .C(\para_9_i_0[27] ), 
        .Y(N_139));
    NOR3 \para_RNO[31]  (.A(N_354), .B(N_353), .C(\para_9_i_0[31] ), 
        .Y(N_128));
    NOR3 \para_RNO_3[16]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[16]_net_1 ), .Y(N_509));
    NOR3A \para_RNO_0[16]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[17]_net_1 ), .Y(N_508));
    NOR3 \para_RNO[12]  (.A(N_364), .B(N_363), .C(\para_9_i_0[12] ), 
        .Y(N_133));
    NOR3 \para_RNO[8]  (.A(N_492), .B(N_491), .C(\para_9_i_0[8] ), .Y(
        N_149));
    OR2A para_reg_18_e (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_540));
    DFN1E0 \para_reg[9]  (.D(dds_configdata[8]), .CLK(GLA), .E(N_540), 
        .Q(\para_reg[9]_net_1 ));
    NOR2B \cs_RNO[6]  (.A(\cs[5]_net_1 ), .B(N_238), .Y(\cs_RNO_0[6] ));
    NOR2 \para_RNO_1[4]  (.A(\para[4]_net_1 ), .B(N_572_1), .Y(N_484));
    NOR2 \para_RNO_1[11]  (.A(\para[11]_net_1 ), .B(N_572_1), .Y(N_503)
        );
    AO1D \para_RNO_2[16]  (.A(dds_configdata[15]), .B(N_540_0), .C(
        N_509), .Y(\para_9_i_0[16] ));
    DFN1E0 \para[29]  (.D(N_143), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[29]_net_1 ));
    OR3 data_RNO_0 (.A(N_239), .B(\cs[4]_net_1 ), .C(\cs[5]_net_1 ), 
        .Y(N_466));
    DFN1 fq_ud (.D(fq_ud_RNO_net_1), .CLK(GLA), .Q(ddsfqud_c));
    NOR2 \para_RNO_1[26]  (.A(\para[26]_net_1 ), .B(N_540_1), .Y(N_523)
        );
    NOR2 \para_RNO_1[17]  (.A(\para[17]_net_1 ), .B(N_540_1), .Y(N_341)
        );
    AO1B state_over_RNO (.A(dds_state_0_state_over), .B(N_539), .C(
        N_238), .Y(state_over_RNO_net_1));
    NOR3 \para_RNO_3[13]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[13]_net_1 ), .Y(N_369));
    NOR3A \para_RNO_0[13]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[14]_net_1 ), .Y(N_368));
    DFN1E0 \para[2]  (.D(N_44), .CLK(GLA), .E(para_1_sqmuxa_1), .Q(
        \para[2]_net_1 ));
    NOR3A \para_RNO_0[22]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[23]_net_1 ), .Y(N_451));
    OR2B para_reg_34_e_0 (.A(top_code_0_dds_load), .B(
        top_code_0_dds_choice), .Y(N_572_0));
    NOR3 \para_RNO_3[15]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para_reg[15]_net_1 ), .Y(N_440));
    NOR2 \para_RNO_1[14]  (.A(\para[14]_net_1 ), .B(N_572_1), .Y(N_371)
        );
    NOR3A \para_RNO_0[15]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[16]_net_1 ), .Y(N_439));
    AO1D \para_RNO_2[13]  (.A(dds_configdata[12]), .B(N_540_0), .C(
        N_369), .Y(\para_9_i_0[13] ));
    NOR3A \para_RNO_0[32]  (.A(i_RNIV2B7[0]), .B(top_code_0_dds_load), 
        .C(\para[33]_net_1 ), .Y(N_528));
    NOR3 \para_RNO[9]  (.A(N_496), .B(N_495), .C(\para_9_i_0[9] ), .Y(
        N_151));
    AO1D \para_RNO_2[15]  (.A(dds_configdata[14]), .B(N_540_0), .C(
        N_440), .Y(\para_9_i_0[15] ));
    AO1D \para_RNO_2[5]  (.A(dds_configdata[4]), .B(N_540_0), .C(N_405)
        , .Y(\para_9_i_0[5] ));
    NOR2 \para_RNO_1[23]  (.A(\para[23]_net_1 ), .B(N_540_1), .Y(N_511)
        );
    NOR3 \para_RNO[15]  (.A(N_439), .B(N_438), .C(\para_9_i_0[15] ), 
        .Y(N_7));
    NOR2 \para_RNO_1[25]  (.A(\para[25]_net_1 ), .B(N_540_1), .Y(N_519)
        );
    
endmodule


module dds_coder(
       i_2,
       count_2,
       count_0,
       i_RNIV2B7,
       GLA,
       dds_change_0_dds_conf,
       dds_change_0_dds_rst
    );
output [3:1] i_2;
input  [4:0] count_2;
input  [7:5] count_0;
output [0:0] i_RNIV2B7;
input  GLA;
input  dds_change_0_dds_conf;
input  dds_change_0_dds_rst;

    wire \i[0]_net_1 , \i_0_0_a2_2[3] , \i_0_0_a2_1[3] , 
        \i_0_0_a2_0_0[1]_net_1 , \i_0_0_a2_4_0[1]_net_1 , N_20, 
        \i_RNO_0[3]_net_1 , \i_RNO_0[2] , N_8_4, N_4, \i_RNO_0[1] , 
        GND, VCC, GND_0, VCC_0;
    
    CLKINT \i_RNIV2B7[0]  (.A(\i[0]_net_1 ), .Y(i_RNIV2B7[0]));
    OR2 \i_0_0_a2_0_0[1]  (.A(count_2[4]), .B(count_0[7]), .Y(
        \i_0_0_a2_0_0[1]_net_1 ));
    DFN1 \i[3]  (.D(\i_RNO_0[3]_net_1 ), .CLK(GLA), .Q(i_2[3]));
    OR3A \i_0_0_a2_4[1]  (.A(\i_0_0_a2_4_0[1]_net_1 ), .B(count_0[6]), 
        .C(count_0[5]), .Y(N_8_4));
    NOR2 \i_RNO_1[3]  (.A(count_2[1]), .B(count_2[3]), .Y(
        \i_0_0_a2_1[3] ));
    DFN1 \i[0]  (.D(N_4), .CLK(GLA), .Q(\i[0]_net_1 ));
    GND GND_i_0 (.Y(GND_0));
    DFN1 \i[2]  (.D(\i_RNO_0[2] ), .CLK(GLA), .Q(i_2[2]));
    VCC VCC_i (.Y(VCC));
    NOR2B \i_RNO[0]  (.A(dds_change_0_dds_rst), .B(
        dds_change_0_dds_conf), .Y(N_4));
    NOR2B \i_0_0_a2_4_0[1]  (.A(count_2[1]), .B(count_2[3]), .Y(
        \i_0_0_a2_4_0[1]_net_1 ));
    NOR3A \i_RNO[3]  (.A(\i_0_0_a2_2[3] ), .B(N_20), .C(count_2[2]), 
        .Y(\i_RNO_0[3]_net_1 ));
    NOR3 \i_RNO[1]  (.A(N_20), .B(count_2[2]), .C(N_8_4), .Y(
        \i_RNO_0[1] ));
    NOR3C \i_RNO_0[3]  (.A(count_0[6]), .B(count_0[5]), .C(
        \i_0_0_a2_1[3] ), .Y(\i_0_0_a2_2[3] ));
    GND GND_i (.Y(GND));
    DFN1 \i[1]  (.D(\i_RNO_0[1] ), .CLK(GLA), .Q(i_2[1]));
    VCC VCC_i_0 (.Y(VCC_0));
    OR3A \i_0_0_a2_0[1]  (.A(dds_change_0_dds_rst), .B(count_2[0]), .C(
        \i_0_0_a2_0_0[1]_net_1 ), .Y(N_20));
    NOR3A \i_RNO[2]  (.A(count_2[2]), .B(N_8_4), .C(N_20), .Y(
        \i_RNO_0[2] ));
    
endmodule


module DDS(
       dds_configdata,
       top_code_0_dds_load,
       top_code_0_dds_choice,
       ddswclk_c,
       ddsfqud_c,
       ddsdata_c,
       ddsreset_c,
       dds_change_0_dds_conf,
       dds_change_0_dds_rst,
       GLA
    );
input  [15:0] dds_configdata;
input  top_code_0_dds_load;
input  top_code_0_dds_choice;
output ddswclk_c;
output ddsfqud_c;
output ddsdata_c;
output ddsreset_c;
input  dds_change_0_dds_conf;
input  dds_change_0_dds_rst;
input  GLA;

    wire \count_2[0] , \count_2[1] , \count_2[2] , \count_2[3] , 
        \count_2[4] , \count_0[5] , \count_0[6] , \count_0[7] , 
        dds_state_0_state_over, \i_2[1] , \i_2[2] , \i_2[3] , 
        \i_RNIV2B7[0] , GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    dds_timer dds_timer_0 (.count_2({\count_2[4] , \count_2[3] , 
        \count_2[2] , \count_2[1] , \count_2[0] }), .count_0({
        \count_0[7] , \count_0[6] , \count_0[5] }), .GLA(GLA), 
        .dds_change_0_dds_rst(dds_change_0_dds_rst), 
        .dds_change_0_dds_conf(dds_change_0_dds_conf), 
        .dds_state_0_state_over(dds_state_0_state_over));
    dds_state dds_state_0 (.i_2({\i_2[3] , \i_2[2] , \i_2[1] }), 
        .dds_configdata({dds_configdata[15], dds_configdata[14], 
        dds_configdata[13], dds_configdata[12], dds_configdata[11], 
        dds_configdata[10], dds_configdata[9], dds_configdata[8], 
        dds_configdata[7], dds_configdata[6], dds_configdata[5], 
        dds_configdata[4], dds_configdata[3], dds_configdata[2], 
        dds_configdata[1], dds_configdata[0]}), .i_RNIV2B7({
        \i_RNIV2B7[0] }), .ddsreset_c(ddsreset_c), .ddsdata_c(
        ddsdata_c), .ddsfqud_c(ddsfqud_c), .ddswclk_c(ddswclk_c), .GLA(
        GLA), .dds_change_0_dds_rst(dds_change_0_dds_rst), 
        .dds_state_0_state_over(dds_state_0_state_over), 
        .top_code_0_dds_choice(top_code_0_dds_choice), 
        .top_code_0_dds_load(top_code_0_dds_load));
    dds_coder dds_coder_0 (.i_2({\i_2[3] , \i_2[2] , \i_2[1] }), 
        .count_2({\count_2[4] , \count_2[3] , \count_2[2] , 
        \count_2[1] , \count_2[0] }), .count_0({\count_0[7] , 
        \count_0[6] , \count_0[5] }), .i_RNIV2B7({\i_RNIV2B7[0] }), 
        .GLA(GLA), .dds_change_0_dds_conf(dds_change_0_dds_conf), 
        .dds_change_0_dds_rst(dds_change_0_dds_rst));
    GND GND_i (.Y(GND));
    
endmodule


module Timer_Cmp(
       dataout,
       timedata,
       cmp_result
    );
input  [21:0] dataout;
input  [21:0] timedata;
output cmp_result;

    wire AO1C_4_Y, AO1C_10_Y, XNOR2_7_Y, NAND3A_0_Y, OR2A_7_Y, 
        AND3_4_Y, XNOR2_19_Y, XNOR2_23_Y, XNOR2_2_Y, XNOR2_21_Y, 
        NOR3A_3_Y, OR2A_2_Y, AO1C_1_Y, OR2A_6_Y, AO1_0_Y, AND3_7_Y, 
        NAND3A_2_Y, NAND3A_6_Y, OR2A_5_Y, AO1C_2_Y, XNOR2_0_Y, 
        AO1C_7_Y, XNOR2_11_Y, OR2A_0_Y, AO1C_8_Y, AO1C_0_Y, OR2A_4_Y, 
        OR2A_11_Y, OR2A_8_Y, NAND3A_7_Y, NOR3A_5_Y, AO1C_3_Y, 
        XNOR2_27_Y, AND3_1_Y, AND3_0_Y, AND3_6_Y, AND3_3_Y, XNOR2_24_Y, 
        XNOR2_20_Y, NOR2A_0_Y, XNOR2_17_Y, NAND3A_5_Y, NOR3A_4_Y, 
        NAND3A_4_Y, XNOR2_25_Y, XNOR2_26_Y, OR2A_13_Y, AO1_2_Y, 
        AND3_5_Y, AO1_4_Y, XNOR2_13_Y, AO1C_9_Y, XNOR2_14_Y, 
        NAND3A_3_Y, NAND3A_10_Y, NOR3A_0_Y, OR2A_12_Y, XNOR2_10_Y, 
        XNOR2_6_Y, AO1_3_Y, NAND3A_1_Y, NAND3A_8_Y, XNOR2_15_Y, 
        XNOR2_16_Y, XNOR2_5_Y, XNOR2_8_Y, OR2A_10_Y, XNOR2_1_Y, 
        AND2_0_Y, AO1_1_Y, XNOR2_28_Y, XNOR2_4_Y, OR2A_3_Y, AND3_8_Y, 
        XNOR2_22_Y, OR2A_9_Y, AO1C_5_Y, XNOR2_9_Y, XNOR2_18_Y, 
        AND2_1_Y, AND3_9_Y, XNOR2_12_Y, AO1C_6_Y, NAND3A_11_Y, 
        AND2_2_Y, AO1D_0_Y, NAND3A_9_Y, AND3_2_Y, NOR3A_2_Y, XNOR2_3_Y, 
        NOR3A_1_Y, OR2A_1_Y, GND, VCC, GND_0, VCC_0;
    
    OR2A OR2A_1 (.A(timedata[8]), .B(dataout[8]), .Y(OR2A_1_Y));
    XNOR2 XNOR2_3 (.A(dataout[3]), .B(timedata[3]), .Y(XNOR2_3_Y));
    OR2A OR2A_10 (.A(dataout[5]), .B(timedata[5]), .Y(OR2A_10_Y));
    AND3 AND3_5 (.A(XNOR2_8_Y), .B(AND3_8_Y), .C(AND2_2_Y), .Y(
        AND3_5_Y));
    NAND3A NAND3A_2 (.A(NOR3A_1_Y), .B(OR2A_1_Y), .C(NAND3A_3_Y), .Y(
        NAND3A_2_Y));
    NAND3A NAND3A_6 (.A(NOR3A_0_Y), .B(OR2A_13_Y), .C(NAND3A_11_Y), .Y(
        NAND3A_6_Y));
    NOR3A NOR3A_1 (.A(OR2A_5_Y), .B(AO1C_7_Y), .C(dataout[6]), .Y(
        NOR3A_1_Y));
    AND3 AND3_2 (.A(XNOR2_3_Y), .B(XNOR2_10_Y), .C(XNOR2_18_Y), .Y(
        AND3_2_Y));
    AO1C AO1C_3 (.A(timedata[13]), .B(dataout[13]), .C(timedata[12]), 
        .Y(AO1C_3_Y));
    AND2 AND2_0 (.A(AND3_1_Y), .B(XNOR2_25_Y), .Y(AND2_0_Y));
    XNOR2 XNOR2_12 (.A(dataout[13]), .B(timedata[13]), .Y(XNOR2_12_Y));
    NOR3A NOR3A_2 (.A(OR2A_7_Y), .B(AO1C_6_Y), .C(dataout[15]), .Y(
        NOR3A_2_Y));
    VCC VCC_i (.Y(VCC));
    NAND3A NAND3A_8 (.A(NOR3A_2_Y), .B(OR2A_11_Y), .C(NAND3A_0_Y), .Y(
        NAND3A_8_Y));
    AO1 AO1_1 (.A(AND2_1_Y), .B(AO1_3_Y), .C(AO1D_0_Y), .Y(AO1_1_Y));
    AND3 AND3_9 (.A(XNOR2_7_Y), .B(XNOR2_4_Y), .C(XNOR2_26_Y), .Y(
        AND3_9_Y));
    XNOR2 XNOR2_22 (.A(dataout[8]), .B(timedata[8]), .Y(XNOR2_22_Y));
    AO1 AO1_4 (.A(AND3_2_Y), .B(NAND3A_9_Y), .C(NAND3A_5_Y), .Y(
        AO1_4_Y));
    NAND3A NAND3A_9 (.A(NOR3A_3_Y), .B(OR2A_4_Y), .C(NAND3A_10_Y), .Y(
        NAND3A_9_Y));
    AO1D AO1D_0 (.A(AO1C_4_Y), .B(AO1C_5_Y), .C(AO1C_8_Y), .Y(AO1D_0_Y)
        );
    AND2 AND2_2 (.A(XNOR2_27_Y), .B(XNOR2_13_Y), .Y(AND2_2_Y));
    NAND3A NAND3A_4 (.A(dataout[4]), .B(timedata[4]), .C(OR2A_10_Y), 
        .Y(NAND3A_4_Y));
    NAND3A NAND3A_11 (.A(dataout[10]), .B(timedata[10]), .C(OR2A_12_Y), 
        .Y(NAND3A_11_Y));
    AO1C AO1C_6 (.A(timedata[16]), .B(dataout[16]), .C(timedata[15]), 
        .Y(AO1C_6_Y));
    AND3 AND3_7 (.A(XNOR2_0_Y), .B(XNOR2_6_Y), .C(XNOR2_16_Y), .Y(
        AND3_7_Y));
    AND3 AND3_6 (.A(XNOR2_24_Y), .B(XNOR2_12_Y), .C(XNOR2_9_Y), .Y(
        AND3_6_Y));
    AND2 AND2_1 (.A(AND3_9_Y), .B(XNOR2_15_Y), .Y(AND2_1_Y));
    XNOR2 XNOR2_9 (.A(dataout[14]), .B(timedata[14]), .Y(XNOR2_9_Y));
    XNOR2 XNOR2_18 (.A(dataout[5]), .B(timedata[5]), .Y(XNOR2_18_Y));
    OR2A OR2A_12 (.A(dataout[11]), .B(timedata[11]), .Y(OR2A_12_Y));
    AO1C AO1C_5 (.A(timedata[20]), .B(dataout[20]), .C(OR2A_9_Y), .Y(
        AO1C_5_Y));
    OR2A OR2A_9 (.A(dataout[19]), .B(timedata[19]), .Y(OR2A_9_Y));
    NAND3A NAND3A_1 (.A(NOR3A_5_Y), .B(OR2A_3_Y), .C(NAND3A_7_Y), .Y(
        NAND3A_1_Y));
    AND3 AND3_0 (.A(XNOR2_14_Y), .B(XNOR2_20_Y), .C(XNOR2_5_Y), .Y(
        AND3_0_Y));
    AND3 AND3_8 (.A(XNOR2_1_Y), .B(XNOR2_28_Y), .C(XNOR2_22_Y), .Y(
        AND3_8_Y));
    OR2A OR2A_3 (.A(timedata[14]), .B(dataout[14]), .Y(OR2A_3_Y));
    XNOR2 XNOR2_4 (.A(dataout[19]), .B(timedata[19]), .Y(XNOR2_4_Y));
    OR2A OR2A_6 (.A(timedata[19]), .B(dataout[19]), .Y(OR2A_6_Y));
    AO1C AO1C_0 (.A(timedata[21]), .B(dataout[21]), .C(NOR2A_0_Y), .Y(
        AO1C_0_Y));
    XNOR2 XNOR2_28 (.A(dataout[7]), .B(timedata[7]), .Y(XNOR2_28_Y));
    AO1 AO1_AGB (.A(AND2_0_Y), .B(AO1_2_Y), .C(AO1_1_Y), .Y(cmp_result)
        );
    XNOR2 XNOR2_1 (.A(dataout[6]), .B(timedata[6]), .Y(XNOR2_1_Y));
    XNOR2 XNOR2_8 (.A(dataout[9]), .B(timedata[9]), .Y(XNOR2_8_Y));
    NOR3A NOR3A_4 (.A(OR2A_10_Y), .B(AO1C_9_Y), .C(dataout[3]), .Y(
        NOR3A_4_Y));
    XNOR2 XNOR2_5 (.A(dataout[20]), .B(timedata[20]), .Y(XNOR2_5_Y));
    XNOR2 XNOR2_16 (.A(dataout[11]), .B(timedata[11]), .Y(XNOR2_16_Y));
    XNOR2 XNOR2_15 (.A(dataout[21]), .B(timedata[21]), .Y(XNOR2_15_Y));
    OR2A OR2A_7 (.A(dataout[17]), .B(timedata[17]), .Y(OR2A_7_Y));
    AO1 AO1_3 (.A(AND3_4_Y), .B(NAND3A_1_Y), .C(NAND3A_8_Y), .Y(
        AO1_3_Y));
    XNOR2 XNOR2_6 (.A(dataout[10]), .B(timedata[10]), .Y(XNOR2_6_Y));
    GND GND_i (.Y(GND));
    XNOR2 XNOR2_10 (.A(dataout[4]), .B(timedata[4]), .Y(XNOR2_10_Y));
    NOR3A NOR3A_0 (.A(OR2A_12_Y), .B(AO1C_2_Y), .C(dataout[9]), .Y(
        NOR3A_0_Y));
    NAND3A NAND3A_10 (.A(dataout[1]), .B(timedata[1]), .C(OR2A_2_Y), 
        .Y(NAND3A_10_Y));
    XNOR2 XNOR2_14 (.A(dataout[18]), .B(timedata[18]), .Y(XNOR2_14_Y));
    NAND3A NAND3A_3 (.A(dataout[7]), .B(timedata[7]), .C(OR2A_5_Y), .Y(
        NAND3A_3_Y));
    XNOR2 XNOR2_2 (.A(dataout[17]), .B(timedata[17]), .Y(XNOR2_2_Y));
    XNOR2 XNOR2_17 (.A(dataout[17]), .B(timedata[17]), .Y(XNOR2_17_Y));
    XNOR2 XNOR2_13 (.A(dataout[11]), .B(timedata[11]), .Y(XNOR2_13_Y));
    AO1 AO1_2 (.A(AND3_5_Y), .B(AO1_4_Y), .C(AO1_0_Y), .Y(AO1_2_Y));
    AO1C AO1C_9 (.A(timedata[4]), .B(dataout[4]), .C(timedata[3]), .Y(
        AO1C_9_Y));
    XNOR2 XNOR2_26 (.A(dataout[20]), .B(timedata[20]), .Y(XNOR2_26_Y));
    XNOR2 XNOR2_25 (.A(dataout[21]), .B(timedata[21]), .Y(XNOR2_25_Y));
    OR2A OR2A_13 (.A(timedata[11]), .B(dataout[11]), .Y(OR2A_13_Y));
    NAND3A NAND3A_5 (.A(NOR3A_4_Y), .B(OR2A_0_Y), .C(NAND3A_4_Y), .Y(
        NAND3A_5_Y));
    AND3 AND3_3 (.A(XNOR2_21_Y), .B(XNOR2_11_Y), .C(XNOR2_17_Y), .Y(
        AND3_3_Y));
    XNOR2 XNOR2_20 (.A(dataout[19]), .B(timedata[19]), .Y(XNOR2_20_Y));
    NOR2A NOR2A_0 (.A(timedata[20]), .B(dataout[20]), .Y(NOR2A_0_Y));
    XNOR2 XNOR2_19 (.A(dataout[15]), .B(timedata[15]), .Y(XNOR2_19_Y));
    XNOR2 XNOR2_24 (.A(dataout[12]), .B(timedata[12]), .Y(XNOR2_24_Y));
    AND3 AND3_1 (.A(AND3_0_Y), .B(AND3_6_Y), .C(AND3_3_Y), .Y(AND3_1_Y)
        );
    XNOR2 XNOR2_27 (.A(dataout[10]), .B(timedata[10]), .Y(XNOR2_27_Y));
    NOR3A NOR3A_5 (.A(OR2A_8_Y), .B(AO1C_3_Y), .C(dataout[12]), .Y(
        NOR3A_5_Y));
    XNOR2 XNOR2_23 (.A(dataout[16]), .B(timedata[16]), .Y(XNOR2_23_Y));
    OR2A OR2A_8 (.A(dataout[14]), .B(timedata[14]), .Y(OR2A_8_Y));
    NAND3A NAND3A_7 (.A(dataout[13]), .B(timedata[13]), .C(OR2A_8_Y), 
        .Y(NAND3A_7_Y));
    OR2A OR2A_11 (.A(timedata[17]), .B(dataout[17]), .Y(OR2A_11_Y));
    OR2A OR2A_4 (.A(timedata[2]), .B(dataout[2]), .Y(OR2A_4_Y));
    OR2A OR2A_0 (.A(timedata[5]), .B(dataout[5]), .Y(OR2A_0_Y));
    AO1C AO1C_8 (.A(dataout[21]), .B(timedata[21]), .C(AO1C_0_Y), .Y(
        AO1C_8_Y));
    AO1C AO1C_1 (.A(timedata[1]), .B(dataout[1]), .C(timedata[0]), .Y(
        AO1C_1_Y));
    XNOR2 XNOR2_11 (.A(dataout[16]), .B(timedata[16]), .Y(XNOR2_11_Y));
    XNOR2 XNOR2_0 (.A(dataout[9]), .B(timedata[9]), .Y(XNOR2_0_Y));
    OR2A OR2A_2 (.A(dataout[2]), .B(timedata[2]), .Y(OR2A_2_Y));
    AO1C AO1C_7 (.A(timedata[7]), .B(dataout[7]), .C(timedata[6]), .Y(
        AO1C_7_Y));
    AO1C AO1C_2 (.A(timedata[10]), .B(dataout[10]), .C(timedata[9]), 
        .Y(AO1C_2_Y));
    OR2A OR2A_5 (.A(dataout[8]), .B(timedata[8]), .Y(OR2A_5_Y));
    AO1 AO1_0 (.A(AND3_7_Y), .B(NAND3A_2_Y), .C(NAND3A_6_Y), .Y(
        AO1_0_Y));
    NOR3A NOR3A_3 (.A(OR2A_2_Y), .B(AO1C_1_Y), .C(dataout[0]), .Y(
        NOR3A_3_Y));
    AO1C AO1C_10 (.A(dataout[18]), .B(timedata[18]), .C(OR2A_6_Y), .Y(
        AO1C_10_Y));
    XNOR2 XNOR2_21 (.A(dataout[15]), .B(timedata[15]), .Y(XNOR2_21_Y));
    XNOR2 XNOR2_7 (.A(dataout[18]), .B(timedata[18]), .Y(XNOR2_7_Y));
    NAND3A NAND3A_0 (.A(dataout[16]), .B(timedata[16]), .C(OR2A_7_Y), 
        .Y(NAND3A_0_Y));
    AND3 AND3_4 (.A(XNOR2_19_Y), .B(XNOR2_23_Y), .C(XNOR2_2_Y), .Y(
        AND3_4_Y));
    AO1C AO1C_4 (.A(timedata[21]), .B(dataout[21]), .C(AO1C_10_Y), .Y(
        AO1C_4_Y));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module timer(
       dataout,
       GLA,
       net_27,
       timer_0_time_up,
       state_switch_0_state_over_n,
       state_switch_0_state_start
    );
input  [21:0] dataout;
input  GLA;
input  net_27;
output timer_0_time_up;
input  state_switch_0_state_over_n;
input  state_switch_0_state_start;

    wire N_95, \timedata[1]_net_1 , \timedata[0]_net_1 , N_87, 
        \timedata[3]_net_1 , \DWACT_FINC_E[0] , N_64, 
        \timedata[8]_net_1 , \DWACT_FINC_E[4] , N_49, 
        \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , time_up_0_sqmuxa_1, 
        time_up_RNO_net_1, cmp_result, \timedata_4[1] , I_5, 
        \timedata_4[2] , I_9, \timedata_4[3] , I_13, \timedata_4[4] , 
        I_20, \timedata_4[5] , I_24, \timedata_4[6] , I_31, 
        \timedata_4[7] , I_38, \timedata_4[8] , I_45, \timedata_4[9] , 
        I_52, \timedata_4[10] , I_56, \timedata_4[11] , I_66, 
        \timedata_4[12] , I_73, \timedata_4[13] , I_77, 
        \timedata_4[14] , I_84, \timedata_4[15] , I_91, 
        \timedata_4[16] , I_98, \timedata_4[17] , I_105, 
        \timedata_4[18] , I_115, \timedata_4[19] , I_122, 
        \timedata_4[20] , I_129, \timedata_4[21] , I_136, 
        \timedata_4[0] , \timedata[2]_net_1 , \timedata[4]_net_1 , 
        \timedata[5]_net_1 , \timedata[6]_net_1 , \timedata[7]_net_1 , 
        \timedata[9]_net_1 , \timedata[10]_net_1 , 
        \timedata[11]_net_1 , \timedata[12]_net_1 , 
        \timedata[13]_net_1 , \timedata[14]_net_1 , 
        \timedata[15]_net_1 , \timedata[16]_net_1 , 
        \timedata[17]_net_1 , \timedata[18]_net_1 , 
        \timedata[19]_net_1 , \timedata[20]_net_1 , 
        \timedata[21]_net_1 , N_4, \DWACT_FINC_E[28] , 
        \DWACT_FINC_E[13] , \DWACT_FINC_E[15] , N_9, 
        \DWACT_FINC_E[14] , N_14, \DWACT_FINC_E[9] , 
        \DWACT_FINC_E[12] , N_19, \DWACT_FINC_E[10] , 
        \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , N_26, \DWACT_FINC_E[11] , 
        N_31, N_36, N_41, \DWACT_FINC_E[8] , N_46, N_54, N_61, 
        \DWACT_FINC_E[3] , N_69, N_74, N_79, \DWACT_FINC_E[1] , N_84, 
        N_92, GND, VCC, GND_0, VCC_0;
    
    XOR2 un2_timedata_I_5 (.A(\timedata[0]_net_1 ), .B(
        \timedata[1]_net_1 ), .Y(I_5));
    NOR3C \timedata_RNO[9]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_52), .Y(\timedata_4[9] ));
    XOR2 un2_timedata_I_13 (.A(N_92), .B(\timedata[3]_net_1 ), .Y(I_13)
        );
    AND3 un2_timedata_I_97 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\timedata[15]_net_1 ), .Y(N_31));
    AND3 un2_timedata_I_87 (.A(\timedata[12]_net_1 ), .B(
        \timedata[13]_net_1 ), .C(\timedata[14]_net_1 ), .Y(
        \DWACT_FINC_E[9] ));
    DFN1 \timedata[14]  (.D(\timedata_4[14] ), .CLK(GLA), .Q(
        \timedata[14]_net_1 ));
    AND3 un2_timedata_I_128 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[14] ), .Y(N_9));
    NOR3C \timedata_RNO[11]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_66), .Y(\timedata_4[11] ));
    NOR3C \timedata_RNO[15]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_91), .Y(\timedata_4[15] ));
    DFN1 \timedata[18]  (.D(\timedata_4[18] ), .CLK(GLA), .Q(
        \timedata[18]_net_1 ));
    DFN1 \timedata[1]  (.D(\timedata_4[1] ), .CLK(GLA), .Q(
        \timedata[1]_net_1 ));
    AND2 un2_timedata_I_125 (.A(\timedata[18]_net_1 ), .B(
        \timedata[19]_net_1 ), .Y(\DWACT_FINC_E[14] ));
    AND3 un2_timedata_I_16 (.A(\timedata[0]_net_1 ), .B(
        \timedata[1]_net_1 ), .C(\timedata[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    NOR3C \timedata_RNO[2]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_9), .Y(\timedata_4[2] ));
    NOR3C \timedata_RNO[13]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_77), .Y(\timedata_4[13] ));
    DFN1 \timedata[9]  (.D(\timedata_4[9] ), .CLK(GLA), .Q(
        \timedata[9]_net_1 ));
    AND3 un2_timedata_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[1] ), .C(\timedata[5]_net_1 ), .Y(N_79));
    XOR2 un2_timedata_I_24 (.A(N_84), .B(\timedata[5]_net_1 ), .Y(I_24)
        );
    VCC VCC_i (.Y(VCC));
    NOR3C \timedata_RNO[21]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_136), .Y(\timedata_4[21] ));
    NOR2B un2_timedata_I_19 (.A(\timedata[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_87));
    AND3 un2_timedata_I_104 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[11] ), .Y(N_26));
    XOR2 un2_timedata_I_77 (.A(N_46), .B(\timedata[13]_net_1 ), .Y(
        I_77));
    AND3 un2_timedata_I_65 (.A(\DWACT_FINC_E[6] ), .B(
        \timedata[9]_net_1 ), .C(\timedata[10]_net_1 ), .Y(N_54));
    XOR2 un2_timedata_I_98 (.A(N_31), .B(\timedata[16]_net_1 ), .Y(
        I_98));
    XOR2 un2_timedata_I_66 (.A(N_54), .B(\timedata[11]_net_1 ), .Y(
        I_66));
    AND3 un2_timedata_I_55 (.A(\DWACT_FINC_E[4] ), .B(
        \timedata[8]_net_1 ), .C(\timedata[9]_net_1 ), .Y(N_61));
    XOR2 un2_timedata_I_45 (.A(N_69), .B(\timedata[8]_net_1 ), .Y(I_45)
        );
    XOR2 un2_timedata_I_9 (.A(N_95), .B(\timedata[2]_net_1 ), .Y(I_9));
    NOR2B un2_timedata_I_8 (.A(\timedata[1]_net_1 ), .B(
        \timedata[0]_net_1 ), .Y(N_95));
    XOR2 un2_timedata_I_56 (.A(N_61), .B(\timedata[10]_net_1 ), .Y(
        I_56));
    AND2 un2_timedata_I_101 (.A(\timedata[15]_net_1 ), .B(
        \timedata[16]_net_1 ), .Y(\DWACT_FINC_E[11] ));
    Timer_Cmp Timer_Cmp_0 (.dataout({dataout[21], dataout[20], 
        dataout[19], dataout[18], dataout[17], dataout[16], 
        dataout[15], dataout[14], dataout[13], dataout[12], 
        dataout[11], dataout[10], dataout[9], dataout[8], dataout[7], 
        dataout[6], dataout[5], dataout[4], dataout[3], dataout[2], 
        dataout[1], dataout[0]}), .timedata({\timedata[21]_net_1 , 
        \timedata[20]_net_1 , \timedata[19]_net_1 , 
        \timedata[18]_net_1 , \timedata[17]_net_1 , 
        \timedata[16]_net_1 , \timedata[15]_net_1 , 
        \timedata[14]_net_1 , \timedata[13]_net_1 , 
        \timedata[12]_net_1 , \timedata[11]_net_1 , 
        \timedata[10]_net_1 , \timedata[9]_net_1 , \timedata[8]_net_1 , 
        \timedata[7]_net_1 , \timedata[6]_net_1 , \timedata[5]_net_1 , 
        \timedata[4]_net_1 , \timedata[3]_net_1 , \timedata[2]_net_1 , 
        \timedata[1]_net_1 , \timedata[0]_net_1 }), .cmp_result(
        cmp_result));
    NOR2B un2_timedata_I_72 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_49));
    AND3 un2_timedata_I_69 (.A(\timedata[9]_net_1 ), .B(
        \timedata[10]_net_1 ), .C(\timedata[11]_net_1 ), .Y(
        \DWACT_FINC_E[7] ));
    NOR3C \timedata_RNO[14]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_84), .Y(\timedata_4[14] ));
    AND3 un2_timedata_I_59 (.A(\timedata[6]_net_1 ), .B(
        \timedata[7]_net_1 ), .C(\timedata[8]_net_1 ), .Y(
        \DWACT_FINC_E[5] ));
    NOR3C \timedata_RNO[6]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_31), .Y(\timedata_4[6] ));
    DFN1 \timedata[8]  (.D(\timedata_4[8] ), .CLK(GLA), .Q(
        \timedata[8]_net_1 ));
    NOR3C \timedata_RNO[10]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_56), .Y(\timedata_4[10] ));
    DFN1 \timedata[17]  (.D(\timedata_4[17] ), .CLK(GLA), .Q(
        \timedata[17]_net_1 ));
    AND3 un2_timedata_I_83 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[8] ), .Y(N_41));
    AND3 un2_timedata_I_34 (.A(\timedata[3]_net_1 ), .B(
        \timedata[4]_net_1 ), .C(\timedata[5]_net_1 ), .Y(
        \DWACT_FINC_E[2] ));
    NOR3C \timedata_RNO[5]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_24), .Y(\timedata_4[5] ));
    NOR3C \timedata_RNO[12]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_73), .Y(\timedata_4[12] ));
    DFN1 \timedata[3]  (.D(\timedata_4[3] ), .CLK(GLA), .Q(
        \timedata[3]_net_1 ));
    AND3 un2_timedata_I_135 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\DWACT_FINC_E[15] ), .Y(N_4));
    XOR2 un2_timedata_I_129 (.A(N_9), .B(\timedata[20]_net_1 ), .Y(
        I_129));
    AND3 un2_timedata_I_44 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_69));
    AND2 un2_timedata_I_27 (.A(\timedata[3]_net_1 ), .B(
        \timedata[4]_net_1 ), .Y(\DWACT_FINC_E[1] ));
    AND3 un2_timedata_I_108 (.A(\timedata[15]_net_1 ), .B(
        \timedata[16]_net_1 ), .C(\timedata[17]_net_1 ), .Y(
        \DWACT_FINC_E[12] ));
    NOR3C \timedata_RNO[20]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_129), .Y(\timedata_4[20] ));
    DFN1 \timedata[16]  (.D(\timedata_4[16] ), .CLK(GLA), .Q(
        \timedata[16]_net_1 ));
    XOR2 un2_timedata_I_31 (.A(N_79), .B(\timedata[6]_net_1 ), .Y(I_31)
        );
    GND GND_i (.Y(GND));
    AND3 un2_timedata_I_90 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\DWACT_FINC_E[9] ), .Y(N_36));
    AND2 un2_timedata_I_80 (.A(\timedata[12]_net_1 ), .B(
        \timedata[13]_net_1 ), .Y(\DWACT_FINC_E[8] ));
    AND3 un2_timedata_I_114 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[10] ), .C(\DWACT_FINC_E[12] ), .Y(N_19));
    DFN1 \timedata[19]  (.D(\timedata_4[19] ), .CLK(GLA), .Q(
        \timedata[19]_net_1 ));
    NOR2B un2_timedata_I_51 (.A(\timedata[8]_net_1 ), .B(
        \DWACT_FINC_E[4] ), .Y(N_64));
    AND2 un2_timedata_I_41 (.A(\timedata[6]_net_1 ), .B(
        \timedata[7]_net_1 ), .Y(\DWACT_FINC_E[3] ));
    XOR2 un2_timedata_I_105 (.A(N_26), .B(\timedata[17]_net_1 ), .Y(
        I_105));
    XOR2 un2_timedata_I_73 (.A(N_49), .B(\timedata[12]_net_1 ), .Y(
        I_73));
    AND3 un2_timedata_I_111 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[28] ));
    NOR3C \timedata_RNO[16]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_98), .Y(\timedata_4[16] ));
    OR3C \timedata_RNO[0]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        \timedata[0]_net_1 ), .Y(\timedata_4[0] ));
    DFN1 \timedata[13]  (.D(\timedata_4[13] ), .CLK(GLA), .Q(
        \timedata[13]_net_1 ));
    NOR3C time_up_RNO (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        cmp_result), .Y(time_up_RNO_net_1));
    NOR3B time_up_RNI6K75 (.A(state_switch_0_state_start), .B(
        state_switch_0_state_over_n), .C(timer_0_time_up), .Y(
        time_up_0_sqmuxa_1));
    NOR3C \timedata_RNO[1]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_5), .Y(\timedata_4[1] ));
    NOR3C \timedata_RNO[18]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_115), .Y(\timedata_4[18] ));
    NOR3C \timedata_RNO[4]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_20), .Y(\timedata_4[4] ));
    DFN1 \timedata[11]  (.D(\timedata_4[11] ), .CLK(GLA), .Q(
        \timedata[11]_net_1 ));
    XOR2 un2_timedata_I_122 (.A(N_14), .B(\timedata[19]_net_1 ), .Y(
        I_122));
    DFN1 time_up (.D(time_up_RNO_net_1), .CLK(GLA), .Q(timer_0_time_up)
        );
    DFN1 \timedata[10]  (.D(\timedata_4[10] ), .CLK(GLA), .Q(
        \timedata[10]_net_1 ));
    AND3 un2_timedata_I_37 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\timedata[6]_net_1 ), .Y(N_74));
    NOR3C \timedata_RNO[8]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_45), .Y(\timedata_4[8] ));
    DFN1 \timedata[5]  (.D(\timedata_4[5] ), .CLK(GLA), .Q(
        \timedata[5]_net_1 ));
    AND3 un2_timedata_I_76 (.A(\DWACT_FINC_E[6] ), .B(
        \DWACT_FINC_E[7] ), .C(\timedata[12]_net_1 ), .Y(N_46));
    AND3 un2_timedata_I_12 (.A(\timedata[0]_net_1 ), .B(
        \timedata[1]_net_1 ), .C(\timedata[2]_net_1 ), .Y(N_92));
    NOR3C \timedata_RNO[7]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_38), .Y(\timedata_4[7] ));
    AND2 un2_timedata_I_94 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .Y(\DWACT_FINC_E[10] ));
    XOR2 un2_timedata_I_84 (.A(N_41), .B(\timedata[14]_net_1 ), .Y(
        I_84));
    NOR3C \timedata_RNO[3]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_13), .Y(\timedata_4[3] ));
    DFN1 \timedata[6]  (.D(\timedata_4[6] ), .CLK(GLA), .Q(
        \timedata[6]_net_1 ));
    XOR2 un2_timedata_I_136 (.A(N_4), .B(\timedata[21]_net_1 ), .Y(
        I_136));
    NOR3C \timedata_RNO[19]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_122), .Y(\timedata_4[19] ));
    AND3 un2_timedata_I_118 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[9] ), .C(\DWACT_FINC_E[12] ), .Y(
        \DWACT_FINC_E[13] ));
    DFN1 \timedata[4]  (.D(\timedata_4[4] ), .CLK(GLA), .Q(
        \timedata[4]_net_1 ));
    AND3 un2_timedata_I_62 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    DFN1 \timedata[15]  (.D(\timedata_4[15] ), .CLK(GLA), .Q(
        \timedata[15]_net_1 ));
    XOR2 un2_timedata_I_52 (.A(N_64), .B(\timedata[9]_net_1 ), .Y(I_52)
        );
    XOR2 un2_timedata_I_91 (.A(N_36), .B(\timedata[15]_net_1 ), .Y(
        I_91));
    AND3 un2_timedata_I_23 (.A(\DWACT_FINC_E[0] ), .B(
        \timedata[3]_net_1 ), .C(\timedata[4]_net_1 ), .Y(N_84));
    AND3 un2_timedata_I_121 (.A(\DWACT_FINC_E[28] ), .B(
        \DWACT_FINC_E[13] ), .C(\timedata[18]_net_1 ), .Y(N_14));
    DFN1 \timedata[12]  (.D(\timedata_4[12] ), .CLK(GLA), .Q(
        \timedata[12]_net_1 ));
    DFN1 \timedata[21]  (.D(\timedata_4[21] ), .CLK(GLA), .Q(
        \timedata[21]_net_1 ));
    DFN1 \timedata[0]  (.D(\timedata_4[0] ), .CLK(GLA), .Q(
        \timedata[0]_net_1 ));
    XOR2 un2_timedata_I_115 (.A(N_19), .B(\timedata[18]_net_1 ), .Y(
        I_115));
    DFN1 \timedata[20]  (.D(\timedata_4[20] ), .CLK(GLA), .Q(
        \timedata[20]_net_1 ));
    XOR2 un2_timedata_I_38 (.A(N_74), .B(\timedata[7]_net_1 ), .Y(I_38)
        );
    NOR3C \timedata_RNO[17]  (.A(net_27), .B(time_up_0_sqmuxa_1), .C(
        I_105), .Y(\timedata_4[17] ));
    DFN1 \timedata[7]  (.D(\timedata_4[7] ), .CLK(GLA), .Q(
        \timedata[7]_net_1 ));
    DFN1 \timedata[2]  (.D(\timedata_4[2] ), .CLK(GLA), .Q(
        \timedata[2]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    AND3 un2_timedata_I_48 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    XOR2 un2_timedata_I_20 (.A(N_87), .B(\timedata[4]_net_1 ), .Y(I_20)
        );
    AND3 un2_timedata_I_132 (.A(\timedata[18]_net_1 ), .B(
        \timedata[19]_net_1 ), .C(\timedata[20]_net_1 ), .Y(
        \DWACT_FINC_E[15] ));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module state_switch(
       dataout,
       timecount_1,
       timecount_0,
       timecount,
       timecount_1_1,
       timecount_1_0,
       timer_top_0_clk_en_noise,
       timer_top_0_clk_en_pluse,
       timer_top_0_clk_en_scale,
       timer_top_0_clk_en_scan,
       timer_top_0_clk_en_st1ms,
       state_switch_0_state_over_n,
       state_switch_0_state_start,
       top_code_0_pluse_str,
       scalestate_0_tetw_pluse,
       noisestate_0_state_over_n,
       scanstate_0_state_over_n,
       timer_0_time_up,
       net_27,
       top_code_0_state_1ms_start,
       top_code_0_scale_start,
       top_code_0_noise_start,
       top_code_0_scan_start,
       plusestate_0_state_over_n,
       GLA,
       timer_top_0_clk_en_scale_0
    );
output [21:0] dataout;
input  [15:0] timecount_1;
input  [19:0] timecount_0;
input  [21:0] timecount;
input  [15:0] timecount_1_1;
input  [15:0] timecount_1_0;
output timer_top_0_clk_en_noise;
output timer_top_0_clk_en_pluse;
output timer_top_0_clk_en_scale;
output timer_top_0_clk_en_scan;
output timer_top_0_clk_en_st1ms;
output state_switch_0_state_over_n;
output state_switch_0_state_start;
input  top_code_0_pluse_str;
input  scalestate_0_tetw_pluse;
input  noisestate_0_state_over_n;
input  scanstate_0_state_over_n;
input  timer_0_time_up;
input  net_27;
input  top_code_0_state_1ms_start;
input  top_code_0_scale_start;
input  top_code_0_noise_start;
input  top_code_0_scan_start;
input  plusestate_0_state_over_n;
input  GLA;
output timer_top_0_clk_en_scale_0;

    wire clk_en_scale_0_0_a2_0_a6_net_1, \dataout_0_0_0_1[13] , N_222, 
        N_225, N_226, \dataout_0_0_0_2[8] , N_292, N_187, 
        \dataout_0_0_0_0[8] , N_291, N_185, \dataout_0_0_0_2[10] , 
        N_192, \dataout_0_0_0_0[10] , N_190, \dataout_0_0_0_2[12] , 
        N_197, \dataout_0_0_0_0[12] , N_195, \dataout_0_0_0_2[14] , 
        N_202, \dataout_0_0_0_0[14] , N_200, \dataout_0_0_0_2[15] , 
        N_219, \dataout_0_0_0_0[15] , N_217, \dataout_0_0_0_2[11] , 
        N_229, \dataout_0_0_0_0[11] , N_227, \dataout_0_0_0_2[9] , 
        N_234, \dataout_0_0_0_0[9] , N_232, \dataout_0_0_0_2[7] , 
        N_239, \dataout_0_0_0_0[7] , N_237, \dataout_0_0_0_2[6] , 
        N_244, \dataout_0_0_0_0[6] , N_242, \dataout_0_0_0_2[5] , 
        N_249, \dataout_0_0_0_0[5] , N_247, \dataout_0_0_0_2[4] , 
        N_254, \dataout_0_0_0_0[4] , N_252, \dataout_0_0_0_2[3] , 
        N_259, \dataout_0_0_0_0[3] , N_257, \dataout_0_0_0_1[2] , 
        N_262, N_265, N_266, \dataout_0_0_0_1[1] , N_267, N_270, N_271, 
        \dataout_0_0_0_2[0] , N_274, \dataout_0_0_0_0[0] , N_272, 
        state_over_n_0_i_0, N_215, state_start5_0_0_1, N_286, N_283, 
        state_start5_0_0_a2_3_0_net_1, state_start5_0_0_a2_1_0_net_1, 
        state_start5_0_0_a2_0_net_1, N_279, N_280, N_277, N_290, N_284, 
        state_start5, \dataout_RNO[0]_net_1 , N_276, 
        \dataout_RNO[1]_net_1 , N_269, N_268, \dataout_RNO[2]_net_1 , 
        N_264, N_263, \dataout_RNO[3]_net_1 , N_261, 
        \dataout_RNO[4]_net_1 , N_256, \dataout_RNO[5]_net_1 , N_251, 
        \dataout_RNO[6]_net_1 , N_246, \dataout_RNO[7]_net_1 , N_241, 
        \dataout_RNO[9]_net_1 , N_236, \dataout_RNO[11]_net_1 , N_231, 
        \dataout_RNO[15]_net_1 , N_221, N_30, N_214, N_213, 
        \dataout_RNO[14]_net_1 , N_203, \dataout_RNO[12]_net_1 , N_198, 
        \dataout_RNO[10]_net_1 , N_193, \dataout_RNO[8]_net_1 , N_188, 
        \dataout_RNO[13]_net_1 , N_224, N_223, clk_en_st1ms_RNO_net_1, 
        clk_en_scan_RNO_net_1, clk_en_pluse_RNO_net_1, 
        clk_en_noise_RNO_net_1, \dataout_RNO[20]_net_1 , 
        \dataout_RNO[21]_net_1 , N_206, N_208, N_210, N_212, 
        \dataout_RNO[16]_net_1 , \dataout_RNO[17]_net_1 , 
        \dataout_RNO[18]_net_1 , \dataout_RNO[19]_net_1 , GND, VCC, 
        GND_0, VCC_0;
    
    AOI1B \dataout_RNO_1[14]  (.A(timecount_1_1[14]), .B(N_291), .C(
        N_200), .Y(\dataout_0_0_0_0[14] ));
    OR3C \dataout_RNO[3]  (.A(N_261), .B(\dataout_0_0_0_0[3] ), .C(
        \dataout_0_0_0_2[3] ), .Y(\dataout_RNO[3]_net_1 ));
    DFN1 \dataout[2]  (.D(\dataout_RNO[2]_net_1 ), .CLK(GLA), .Q(
        dataout[2]));
    OR2B \dataout_RNO_0[8]  (.A(timecount[8]), .B(N_283), .Y(N_188));
    OR2B \dataout_RNO_3[14]  (.A(timecount_0[14]), .B(N_286), .Y(N_200)
        );
    AO1B \dataout_RNO[18]  (.A(timecount_0[18]), .B(N_286), .C(N_210), 
        .Y(\dataout_RNO[18]_net_1 ));
    OR2B \dataout_RNO_3[7]  (.A(timecount_0[7]), .B(N_286), .Y(N_237));
    OR2B \dataout_RNO_3[4]  (.A(timecount_0[4]), .B(N_286), .Y(N_252));
    OR2B \dataout_RNO_0[11]  (.A(timecount[11]), .B(N_283), .Y(N_231));
    DFN1 \dataout[1]  (.D(\dataout_RNO[1]_net_1 ), .CLK(GLA), .Q(
        dataout[1]));
    DFN1 \dataout[21]  (.D(\dataout_RNO[21]_net_1 ), .CLK(GLA), .Q(
        dataout[21]));
    OR2B \dataout_RNO_0[4]  (.A(timecount[4]), .B(N_283), .Y(N_256));
    OR2B \dataout_RNO_3[6]  (.A(timecount_0[6]), .B(N_286), .Y(N_242));
    AOI1B \dataout_RNO_2[15]  (.A(timecount_1_0[15]), .B(N_292), .C(
        N_219), .Y(\dataout_0_0_0_2[15] ));
    AOI1B \dataout_RNO_1[4]  (.A(timecount_1_1[4]), .B(N_291), .C(
        N_252), .Y(\dataout_0_0_0_0[4] ));
    OR2B \dataout_RNO_1[2]  (.A(timecount_1_0[2]), .B(N_292), .Y(N_263)
        );
    OR3C \dataout_RNO[4]  (.A(N_256), .B(\dataout_0_0_0_0[4] ), .C(
        \dataout_0_0_0_2[4] ), .Y(\dataout_RNO[4]_net_1 ));
    OR3C \dataout_RNO[0]  (.A(N_276), .B(\dataout_0_0_0_0[0] ), .C(
        \dataout_0_0_0_2[0] ), .Y(\dataout_RNO[0]_net_1 ));
    OR3C \dataout_RNO[2]  (.A(N_264), .B(N_263), .C(
        \dataout_0_0_0_1[2] ), .Y(\dataout_RNO[2]_net_1 ));
    OR2B \dataout_RNO_0[10]  (.A(timecount[10]), .B(N_283), .Y(N_193));
    DFN1 \dataout[0]  (.D(\dataout_RNO[0]_net_1 ), .CLK(GLA), .Q(
        dataout[0]));
    OR2B \dataout_RNO_4[12]  (.A(timecount_1[12]), .B(N_290), .Y(N_197)
        );
    OR3C \dataout_RNO[15]  (.A(N_221), .B(\dataout_0_0_0_0[15] ), .C(
        \dataout_0_0_0_2[15] ), .Y(\dataout_RNO[15]_net_1 ));
    AOI1B \dataout_RNO_1[0]  (.A(timecount_1_1[0]), .B(N_291), .C(
        N_272), .Y(\dataout_0_0_0_0[0] ));
    DFN1 \dataout[14]  (.D(\dataout_RNO[14]_net_1 ), .CLK(GLA), .Q(
        dataout[14]));
    AOI1B \dataout_RNO_2[6]  (.A(timecount_1_0[6]), .B(N_292), .C(
        N_244), .Y(\dataout_0_0_0_2[6] ));
    DFN1 \dataout[3]  (.D(\dataout_RNO[3]_net_1 ), .CLK(GLA), .Q(
        dataout[3]));
    OR3C \dataout_RNO[8]  (.A(N_188), .B(\dataout_0_0_0_0[8] ), .C(
        \dataout_0_0_0_2[8] ), .Y(\dataout_RNO[8]_net_1 ));
    OR2B \dataout_RNO_3[8]  (.A(timecount_0[8]), .B(N_286), .Y(N_185));
    OR2A state_start5_0_0_a2_3_0 (.A(top_code_0_scan_start), .B(
        top_code_0_noise_start), .Y(state_start5_0_0_a2_3_0_net_1));
    OR2B \dataout_RNO_3[3]  (.A(timecount_0[3]), .B(N_286), .Y(N_257));
    OR2B \dataout_RNO_4[8]  (.A(timecount_1[8]), .B(N_290), .Y(N_187));
    OR3C \dataout_RNO[10]  (.A(N_193), .B(\dataout_0_0_0_0[10] ), .C(
        \dataout_0_0_0_2[10] ), .Y(\dataout_RNO[10]_net_1 ));
    AOI1B \dataout_RNO_1[8]  (.A(timecount_1_1[8]), .B(N_291), .C(
        N_185), .Y(\dataout_0_0_0_0[8] ));
    OR2B \dataout_RNO_1[1]  (.A(timecount_1_0[1]), .B(N_292), .Y(N_268)
        );
    OR3A state_start5_0_0_a2_0_0 (.A(top_code_0_scale_start), .B(
        top_code_0_noise_start), .C(top_code_0_scan_start), .Y(
        state_start5_0_0_a2_0_net_1));
    NOR2A state_over_n_RNO_3 (.A(N_283), .B(scalestate_0_tetw_pluse), 
        .Y(N_215));
    NOR2A state_over_n_RNO_1 (.A(N_292), .B(scanstate_0_state_over_n), 
        .Y(N_213));
    DFN1 clk_en_scan (.D(clk_en_scan_RNO_net_1), .CLK(GLA), .Q(
        timer_top_0_clk_en_scan));
    OR2B \dataout_RNO_0[2]  (.A(timecount_1[2]), .B(N_290), .Y(N_264));
    AOI1B \dataout_RNO_2[3]  (.A(timecount_1_0[3]), .B(N_292), .C(
        N_259), .Y(\dataout_0_0_0_2[3] ));
    OR2B \dataout_RNO_0[5]  (.A(timecount[5]), .B(N_283), .Y(N_251));
    AOI1B \dataout_RNO_1[5]  (.A(timecount_1_1[5]), .B(N_291), .C(
        N_247), .Y(\dataout_0_0_0_0[5] ));
    DFN1 clk_en_noise (.D(clk_en_noise_RNO_net_1), .CLK(GLA), .Q(
        timer_top_0_clk_en_noise));
    OR2B \dataout_RNO_0[0]  (.A(timecount[0]), .B(N_283), .Y(N_276));
    DFN1 \dataout[17]  (.D(\dataout_RNO[17]_net_1 ), .CLK(GLA), .Q(
        dataout[17]));
    OR2B \dataout_RNO_0[1]  (.A(timecount_1[1]), .B(N_290), .Y(N_269));
    NOR2A clk_en_pluse_RNO (.A(timer_0_time_up), .B(N_284), .Y(
        clk_en_pluse_RNO_net_1));
    GND GND_i (.Y(GND));
    DFN1 clk_en_pluse (.D(clk_en_pluse_RNO_net_1), .CLK(GLA), .Q(
        timer_top_0_clk_en_pluse));
    NOR3 state_start5_0_0_a2_1 (.A(N_279), .B(top_code_0_scale_start), 
        .C(state_start5_0_0_a2_1_0_net_1), .Y(N_290));
    OR2B \dataout_RNO_3[5]  (.A(timecount_0[5]), .B(N_286), .Y(N_247));
    AOI1B \dataout_RNO_1[12]  (.A(timecount_1_1[12]), .B(N_291), .C(
        N_195), .Y(\dataout_0_0_0_0[12] ));
    NOR3C clk_en_st1ms_RNO (.A(net_27), .B(timer_0_time_up), .C(
        top_code_0_state_1ms_start), .Y(clk_en_st1ms_RNO_net_1));
    OR3C \dataout_RNO[11]  (.A(N_231), .B(\dataout_0_0_0_0[11] ), .C(
        \dataout_0_0_0_2[11] ), .Y(\dataout_RNO[11]_net_1 ));
    OR2B \dataout_RNO_0[18]  (.A(timecount[18]), .B(N_283), .Y(N_210));
    OR2B \dataout_RNO_0[14]  (.A(timecount[14]), .B(N_283), .Y(N_203));
    NOR3A state_start5_0_0_a2_0 (.A(top_code_0_state_1ms_start), .B(
        N_280), .C(N_277), .Y(N_286));
    OR2B \dataout_RNO_4[15]  (.A(timecount_1[15]), .B(N_290), .Y(N_219)
        );
    VCC VCC_i_0 (.Y(VCC_0));
    OR2B \dataout_RNO_3[12]  (.A(timecount_0[12]), .B(N_286), .Y(N_195)
        );
    OR3C \dataout_RNO[9]  (.A(N_236), .B(\dataout_0_0_0_0[9] ), .C(
        \dataout_0_0_0_2[9] ), .Y(\dataout_RNO[9]_net_1 ));
    OR2B \dataout_RNO_3[9]  (.A(timecount_0[9]), .B(N_286), .Y(N_232));
    NOR3C \dataout_RNO_2[1]  (.A(N_267), .B(N_270), .C(N_271), .Y(
        \dataout_0_0_0_1[1] ));
    OR3C \dataout_RNO[6]  (.A(N_246), .B(\dataout_0_0_0_0[6] ), .C(
        \dataout_0_0_0_2[6] ), .Y(\dataout_RNO[6]_net_1 ));
    AOI1B \dataout_RNO_1[3]  (.A(timecount_1_1[3]), .B(N_291), .C(
        N_257), .Y(\dataout_0_0_0_0[3] ));
    AOI1B \dataout_RNO_1[6]  (.A(timecount_1_1[6]), .B(N_291), .C(
        N_242), .Y(\dataout_0_0_0_0[6] ));
    DFN1 \dataout[10]  (.D(\dataout_RNO[10]_net_1 ), .CLK(GLA), .Q(
        dataout[10]));
    DFN1 \dataout[6]  (.D(\dataout_RNO[6]_net_1 ), .CLK(GLA), .Q(
        dataout[6]));
    OR2B \dataout_RNO_3[0]  (.A(timecount_0[0]), .B(N_286), .Y(N_272));
    OR3C \dataout_RNO[13]  (.A(N_224), .B(N_223), .C(
        \dataout_0_0_0_1[13] ), .Y(\dataout_RNO[13]_net_1 ));
    DFN1 state_over_n (.D(N_30), .CLK(GLA), .Q(
        state_switch_0_state_over_n));
    AO1B \dataout_RNO[19]  (.A(timecount_0[19]), .B(N_286), .C(N_212), 
        .Y(\dataout_RNO[19]_net_1 ));
    NOR3C \dataout_RNO_2[13]  (.A(N_222), .B(N_225), .C(N_226), .Y(
        \dataout_0_0_0_1[13] ));
    VCC VCC_i (.Y(VCC));
    OR3A state_start_RNO (.A(state_start5_0_0_1), .B(N_292), .C(N_290), 
        .Y(state_start5));
    OR2B \dataout_RNO_4[2]  (.A(timecount_1_1[2]), .B(N_291), .Y(N_265)
        );
    AOI1B \dataout_RNO_1[15]  (.A(timecount_1_1[15]), .B(N_291), .C(
        N_217), .Y(\dataout_0_0_0_0[15] ));
    DFN1 clk_en_scale (.D(clk_en_scale_0_0_a2_0_a6_net_1), .CLK(GLA), 
        .Q(timer_top_0_clk_en_scale));
    OR2B \dataout_RNO_4[1]  (.A(timecount_1_1[1]), .B(N_291), .Y(N_270)
        );
    AOI1B \dataout_RNO_2[11]  (.A(timecount_1_0[11]), .B(N_292), .C(
        N_229), .Y(\dataout_0_0_0_2[11] ));
    AO1B \dataout_RNO[17]  (.A(timecount_0[17]), .B(N_286), .C(N_208), 
        .Y(\dataout_RNO[17]_net_1 ));
    DFN1 \dataout[5]  (.D(\dataout_RNO[5]_net_1 ), .CLK(GLA), .Q(
        dataout[5]));
    NOR3 state_start5_0_0_a2_3 (.A(N_279), .B(top_code_0_scale_start), 
        .C(state_start5_0_0_a2_3_0_net_1), .Y(N_292));
    OR2B \dataout_RNO_3[15]  (.A(timecount_0[15]), .B(N_286), .Y(N_217)
        );
    OR2B \dataout_RNO_0[9]  (.A(timecount[9]), .B(N_283), .Y(N_236));
    DFN1 \dataout[7]  (.D(\dataout_RNO[7]_net_1 ), .CLK(GLA), .Q(
        dataout[7]));
    NOR3 state_start_RNO_0 (.A(N_286), .B(N_291), .C(N_283), .Y(
        state_start5_0_0_1));
    AOI1B \dataout_RNO_2[10]  (.A(timecount_1_0[10]), .B(N_292), .C(
        N_192), .Y(\dataout_0_0_0_2[10] ));
    OR2B \dataout_RNO_4[7]  (.A(timecount_1[7]), .B(N_290), .Y(N_239));
    OR2B \dataout_RNO_0[19]  (.A(timecount[19]), .B(N_283), .Y(N_212));
    NOR3C clk_en_noise_RNO (.A(net_27), .B(timer_0_time_up), .C(
        top_code_0_noise_start), .Y(clk_en_noise_RNO_net_1));
    AOI1B \dataout_RNO_2[4]  (.A(timecount_1_0[4]), .B(N_292), .C(
        N_254), .Y(\dataout_0_0_0_2[4] ));
    OR2B \dataout_RNO_0[12]  (.A(timecount[12]), .B(N_283), .Y(N_198));
    AOI1B \dataout_RNO_2[7]  (.A(timecount_1_0[7]), .B(N_292), .C(
        N_239), .Y(\dataout_0_0_0_2[7] ));
    OR2B \dataout_RNO_5[1]  (.A(timecount[1]), .B(N_283), .Y(N_271));
    OR2B \dataout_RNO_0[6]  (.A(timecount[6]), .B(N_283), .Y(N_246));
    OR2B \dataout_RNO_4[13]  (.A(timecount_1_1[13]), .B(N_291), .Y(
        N_225));
    NOR2 state_start5_0_0_a2 (.A(state_start5_0_0_a2_0_net_1), .B(
        N_279), .Y(N_283));
    DFN1 \dataout[15]  (.D(\dataout_RNO[15]_net_1 ), .CLK(GLA), .Q(
        dataout[15]));
    AOI1B \dataout_RNO_2[5]  (.A(timecount_1_0[5]), .B(N_292), .C(
        N_249), .Y(\dataout_0_0_0_2[5] ));
    NOR3 state_over_n_RNO (.A(N_214), .B(N_213), .C(state_over_n_0_i_0)
        , .Y(N_30));
    OR2B \dataout_RNO_4[11]  (.A(timecount_1[11]), .B(N_290), .Y(N_229)
        );
    OR2A state_start5_0_0_a2_12 (.A(net_27), .B(top_code_0_pluse_str), 
        .Y(N_277));
    OR2B \dataout_RNO_5[2]  (.A(timecount[2]), .B(N_283), .Y(N_266));
    DFN1 \dataout[4]  (.D(\dataout_RNO[4]_net_1 ), .CLK(GLA), .Q(
        dataout[4]));
    AOI1B \dataout_RNO_2[14]  (.A(timecount_1_0[14]), .B(N_292), .C(
        N_202), .Y(\dataout_0_0_0_2[14] ));
    DFN1 \dataout[11]  (.D(\dataout_RNO[11]_net_1 ), .CLK(GLA), .Q(
        dataout[11]));
    DFN1 \dataout[12]  (.D(\dataout_RNO[12]_net_1 ), .CLK(GLA), .Q(
        dataout[12]));
    GND GND_i_0 (.Y(GND_0));
    OR2B \dataout_RNO_0[15]  (.A(timecount[15]), .B(N_283), .Y(N_221));
    OR2B \dataout_RNO_5[13]  (.A(timecount[13]), .B(N_283), .Y(N_226));
    NOR2A state_over_n_RNO_0 (.A(N_290), .B(noisestate_0_state_over_n), 
        .Y(N_214));
    OR2B \dataout_RNO_0[3]  (.A(timecount[3]), .B(N_283), .Y(N_261));
    AOI1B \dataout_RNO_2[0]  (.A(timecount_1_0[0]), .B(N_292), .C(
        N_274), .Y(\dataout_0_0_0_2[0] ));
    OR2B \dataout_RNO_4[3]  (.A(timecount_1[3]), .B(N_290), .Y(N_259));
    DFN1 \dataout[9]  (.D(\dataout_RNO[9]_net_1 ), .CLK(GLA), .Q(
        dataout[9]));
    OR2B \dataout_RNO_4[10]  (.A(timecount_1[10]), .B(N_290), .Y(N_192)
        );
    OR3A state_start5_0_0_a2_4 (.A(net_27), .B(top_code_0_pluse_str), 
        .C(top_code_0_state_1ms_start), .Y(N_279));
    OR2B \dataout_RNO_4[0]  (.A(timecount_1[0]), .B(N_290), .Y(N_274));
    DFN1 \dataout[13]  (.D(\dataout_RNO[13]_net_1 ), .CLK(GLA), .Q(
        dataout[13]));
    DFN1 \dataout[20]  (.D(\dataout_RNO[20]_net_1 ), .CLK(GLA), .Q(
        dataout[20]));
    AOI1B \dataout_RNO_1[9]  (.A(timecount_1_1[9]), .B(N_291), .C(
        N_232), .Y(\dataout_0_0_0_0[9] ));
    AOI1B \dataout_RNO_2[9]  (.A(timecount_1_0[9]), .B(N_292), .C(
        N_234), .Y(\dataout_0_0_0_2[9] ));
    OR2B \dataout_RNO_1[13]  (.A(timecount_1_0[13]), .B(N_292), .Y(
        N_223));
    DFN1 \dataout[18]  (.D(\dataout_RNO[18]_net_1 ), .CLK(GLA), .Q(
        dataout[18]));
    OR2B \dataout_RNO_3[13]  (.A(timecount_0[13]), .B(N_286), .Y(N_222)
        );
    OR3C \dataout_RNO[5]  (.A(N_251), .B(\dataout_0_0_0_0[5] ), .C(
        \dataout_0_0_0_2[5] ), .Y(\dataout_RNO[5]_net_1 ));
    OR3C \dataout_RNO[14]  (.A(N_203), .B(\dataout_0_0_0_0[14] ), .C(
        \dataout_0_0_0_2[14] ), .Y(\dataout_RNO[14]_net_1 ));
    AOI1B \dataout_RNO_1[11]  (.A(timecount_1_1[11]), .B(N_291), .C(
        N_227), .Y(\dataout_0_0_0_0[11] ));
    OR2B \dataout_RNO_4[5]  (.A(timecount_1[5]), .B(N_290), .Y(N_249));
    OR2B \dataout_RNO_3[11]  (.A(timecount_0[11]), .B(N_286), .Y(N_227)
        );
    OR2B \dataout_RNO_0[7]  (.A(timecount[7]), .B(N_283), .Y(N_241));
    NOR2B \dataout_RNO[20]  (.A(timecount[20]), .B(N_283), .Y(
        \dataout_RNO[20]_net_1 ));
    OR3C \dataout_RNO[1]  (.A(N_269), .B(N_268), .C(
        \dataout_0_0_0_1[1] ), .Y(\dataout_RNO[1]_net_1 ));
    OR3 state_start5_0_0_a2_5 (.A(top_code_0_noise_start), .B(
        top_code_0_scan_start), .C(top_code_0_scale_start), .Y(N_280));
    DFN1 clk_en_scale_0 (.D(clk_en_scale_0_0_a2_0_a6_net_1), .CLK(GLA), 
        .Q(timer_top_0_clk_en_scale_0));
    NOR3 state_start5_0_0_a2_2 (.A(N_280), .B(
        top_code_0_state_1ms_start), .C(N_284), .Y(N_291));
    OR2B \dataout_RNO_0[16]  (.A(timecount[16]), .B(N_283), .Y(N_206));
    AOI1B \dataout_RNO_1[7]  (.A(timecount_1_1[7]), .B(N_291), .C(
        N_237), .Y(\dataout_0_0_0_0[7] ));
    AOI1B \dataout_RNO_1[10]  (.A(timecount_1_1[10]), .B(N_291), .C(
        N_190), .Y(\dataout_0_0_0_0[10] ));
    NOR3C clk_en_scan_RNO (.A(net_27), .B(timer_0_time_up), .C(
        top_code_0_scan_start), .Y(clk_en_scan_RNO_net_1));
    OR2B \dataout_RNO_4[14]  (.A(timecount_1[14]), .B(N_290), .Y(N_202)
        );
    DFN1 \dataout[16]  (.D(\dataout_RNO[16]_net_1 ), .CLK(GLA), .Q(
        dataout[16]));
    OR2B \dataout_RNO_3[10]  (.A(timecount_0[10]), .B(N_286), .Y(N_190)
        );
    OR2B \dataout_RNO_0[17]  (.A(timecount[17]), .B(N_283), .Y(N_208));
    AO1B \dataout_RNO[16]  (.A(timecount_0[16]), .B(N_286), .C(N_206), 
        .Y(\dataout_RNO[16]_net_1 ));
    NOR2B \dataout_RNO[21]  (.A(timecount[21]), .B(N_283), .Y(
        \dataout_RNO[21]_net_1 ));
    DFN1 \dataout[8]  (.D(\dataout_RNO[8]_net_1 ), .CLK(GLA), .Q(
        dataout[8]));
    AOI1B \dataout_RNO_2[12]  (.A(timecount_1_0[12]), .B(N_292), .C(
        N_197), .Y(\dataout_0_0_0_2[12] ));
    OR2A state_start5_0_0_a2_1_0 (.A(top_code_0_noise_start), .B(
        top_code_0_scan_start), .Y(state_start5_0_0_a2_1_0_net_1));
    DFN1 \dataout[19]  (.D(\dataout_RNO[19]_net_1 ), .CLK(GLA), .Q(
        dataout[19]));
    AO1A state_over_n_RNO_2 (.A(plusestate_0_state_over_n), .B(N_291), 
        .C(N_215), .Y(state_over_n_0_i_0));
    NOR3C \dataout_RNO_2[2]  (.A(N_262), .B(N_265), .C(N_266), .Y(
        \dataout_0_0_0_1[2] ));
    OR2B \dataout_RNO_4[6]  (.A(timecount_1[6]), .B(N_290), .Y(N_244));
    OR2B \dataout_RNO_3[1]  (.A(timecount_0[1]), .B(N_286), .Y(N_267));
    OR2B \dataout_RNO_3[2]  (.A(timecount_0[2]), .B(N_286), .Y(N_262));
    NOR3C clk_en_scale_0_0_a2_0_a6 (.A(net_27), .B(timer_0_time_up), 
        .C(top_code_0_scale_start), .Y(clk_en_scale_0_0_a2_0_a6_net_1));
    OR2B \dataout_RNO_4[9]  (.A(timecount_1[9]), .B(N_290), .Y(N_234));
    OR2B \dataout_RNO_4[4]  (.A(timecount_1[4]), .B(N_290), .Y(N_254));
    AOI1B \dataout_RNO_2[8]  (.A(timecount_1_0[8]), .B(N_292), .C(
        N_187), .Y(\dataout_0_0_0_2[8] ));
    DFN1 state_start (.D(state_start5), .CLK(GLA), .Q(
        state_switch_0_state_start));
    OR3C \dataout_RNO[7]  (.A(N_241), .B(\dataout_0_0_0_0[7] ), .C(
        \dataout_0_0_0_2[7] ), .Y(\dataout_RNO[7]_net_1 ));
    OR3C \dataout_RNO[12]  (.A(N_198), .B(\dataout_0_0_0_0[12] ), .C(
        \dataout_0_0_0_2[12] ), .Y(\dataout_RNO[12]_net_1 ));
    OR2B \dataout_RNO_0[13]  (.A(timecount_1[13]), .B(N_290), .Y(N_224)
        );
    DFN1 clk_en_st1ms (.D(clk_en_st1ms_RNO_net_1), .CLK(GLA), .Q(
        timer_top_0_clk_en_st1ms));
    OR2B clk_en_pluse_0_0_a2_0_a2 (.A(top_code_0_pluse_str), .B(net_27)
        , .Y(N_284));
    
endmodule


module timer_top(
       timecount_1_0,
       timecount_1_1,
       timecount,
       timecount_0,
       timecount_1,
       timer_top_0_clk_en_scale_0,
       plusestate_0_state_over_n,
       top_code_0_scan_start,
       top_code_0_noise_start,
       top_code_0_scale_start,
       top_code_0_state_1ms_start,
       scanstate_0_state_over_n,
       noisestate_0_state_over_n,
       scalestate_0_tetw_pluse,
       top_code_0_pluse_str,
       timer_top_0_clk_en_st1ms,
       timer_top_0_clk_en_scan,
       timer_top_0_clk_en_scale,
       timer_top_0_clk_en_pluse,
       timer_top_0_clk_en_noise,
       net_27,
       GLA
    );
input  [15:0] timecount_1_0;
input  [15:0] timecount_1_1;
input  [21:0] timecount;
input  [19:0] timecount_0;
input  [15:0] timecount_1;
output timer_top_0_clk_en_scale_0;
input  plusestate_0_state_over_n;
input  top_code_0_scan_start;
input  top_code_0_noise_start;
input  top_code_0_scale_start;
input  top_code_0_state_1ms_start;
input  scanstate_0_state_over_n;
input  noisestate_0_state_over_n;
input  scalestate_0_tetw_pluse;
input  top_code_0_pluse_str;
output timer_top_0_clk_en_st1ms;
output timer_top_0_clk_en_scan;
output timer_top_0_clk_en_scale;
output timer_top_0_clk_en_pluse;
output timer_top_0_clk_en_noise;
input  net_27;
input  GLA;

    wire \dataout[0] , \dataout[1] , \dataout[2] , \dataout[3] , 
        \dataout[4] , \dataout[5] , \dataout[6] , \dataout[7] , 
        \dataout[8] , \dataout[9] , \dataout[10] , \dataout[11] , 
        \dataout[12] , \dataout[13] , \dataout[14] , \dataout[15] , 
        \dataout[16] , \dataout[17] , \dataout[18] , \dataout[19] , 
        \dataout[20] , \dataout[21] , timer_0_time_up, 
        state_switch_0_state_over_n, state_switch_0_state_start, GND, 
        VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    timer timer_0 (.dataout({\dataout[21] , \dataout[20] , 
        \dataout[19] , \dataout[18] , \dataout[17] , \dataout[16] , 
        \dataout[15] , \dataout[14] , \dataout[13] , \dataout[12] , 
        \dataout[11] , \dataout[10] , \dataout[9] , \dataout[8] , 
        \dataout[7] , \dataout[6] , \dataout[5] , \dataout[4] , 
        \dataout[3] , \dataout[2] , \dataout[1] , \dataout[0] }), .GLA(
        GLA), .net_27(net_27), .timer_0_time_up(timer_0_time_up), 
        .state_switch_0_state_over_n(state_switch_0_state_over_n), 
        .state_switch_0_state_start(state_switch_0_state_start));
    state_switch state_switch_0 (.dataout({\dataout[21] , 
        \dataout[20] , \dataout[19] , \dataout[18] , \dataout[17] , 
        \dataout[16] , \dataout[15] , \dataout[14] , \dataout[13] , 
        \dataout[12] , \dataout[11] , \dataout[10] , \dataout[9] , 
        \dataout[8] , \dataout[7] , \dataout[6] , \dataout[5] , 
        \dataout[4] , \dataout[3] , \dataout[2] , \dataout[1] , 
        \dataout[0] }), .timecount_1({timecount_1[15], timecount_1[14], 
        timecount_1[13], timecount_1[12], timecount_1[11], 
        timecount_1[10], timecount_1[9], timecount_1[8], 
        timecount_1[7], timecount_1[6], timecount_1[5], timecount_1[4], 
        timecount_1[3], timecount_1[2], timecount_1[1], timecount_1[0]})
        , .timecount_0({timecount_0[19], timecount_0[18], 
        timecount_0[17], timecount_0[16], timecount_0[15], 
        timecount_0[14], timecount_0[13], timecount_0[12], 
        timecount_0[11], timecount_0[10], timecount_0[9], 
        timecount_0[8], timecount_0[7], timecount_0[6], timecount_0[5], 
        timecount_0[4], timecount_0[3], timecount_0[2], timecount_0[1], 
        timecount_0[0]}), .timecount({timecount[21], timecount[20], 
        timecount[19], timecount[18], timecount[17], timecount[16], 
        timecount[15], timecount[14], timecount[13], timecount[12], 
        timecount[11], timecount[10], timecount[9], timecount[8], 
        timecount[7], timecount[6], timecount[5], timecount[4], 
        timecount[3], timecount[2], timecount[1], timecount[0]}), 
        .timecount_1_1({timecount_1_1[15], timecount_1_1[14], 
        timecount_1_1[13], timecount_1_1[12], timecount_1_1[11], 
        timecount_1_1[10], timecount_1_1[9], timecount_1_1[8], 
        timecount_1_1[7], timecount_1_1[6], timecount_1_1[5], 
        timecount_1_1[4], timecount_1_1[3], timecount_1_1[2], 
        timecount_1_1[1], timecount_1_1[0]}), .timecount_1_0({
        timecount_1_0[15], timecount_1_0[14], timecount_1_0[13], 
        timecount_1_0[12], timecount_1_0[11], timecount_1_0[10], 
        timecount_1_0[9], timecount_1_0[8], timecount_1_0[7], 
        timecount_1_0[6], timecount_1_0[5], timecount_1_0[4], 
        timecount_1_0[3], timecount_1_0[2], timecount_1_0[1], 
        timecount_1_0[0]}), .timer_top_0_clk_en_noise(
        timer_top_0_clk_en_noise), .timer_top_0_clk_en_pluse(
        timer_top_0_clk_en_pluse), .timer_top_0_clk_en_scale(
        timer_top_0_clk_en_scale), .timer_top_0_clk_en_scan(
        timer_top_0_clk_en_scan), .timer_top_0_clk_en_st1ms(
        timer_top_0_clk_en_st1ms), .state_switch_0_state_over_n(
        state_switch_0_state_over_n), .state_switch_0_state_start(
        state_switch_0_state_start), .top_code_0_pluse_str(
        top_code_0_pluse_str), .scalestate_0_tetw_pluse(
        scalestate_0_tetw_pluse), .noisestate_0_state_over_n(
        noisestate_0_state_over_n), .scanstate_0_state_over_n(
        scanstate_0_state_over_n), .timer_0_time_up(timer_0_time_up), 
        .net_27(net_27), .top_code_0_state_1ms_start(
        top_code_0_state_1ms_start), .top_code_0_scale_start(
        top_code_0_scale_start), .top_code_0_noise_start(
        top_code_0_noise_start), .top_code_0_scan_start(
        top_code_0_scan_start), .plusestate_0_state_over_n(
        plusestate_0_state_over_n), .GLA(GLA), 
        .timer_top_0_clk_en_scale_0(timer_top_0_clk_en_scale_0));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module add_reg_add_reg_2_1(
       addresult_RNI8MQ7,
       addresult_RNIFE5C,
       signal_data_0_iv_i_2,
       addresult_RNIBOIB,
       signal_data_0_iv_i_5,
       signal_data_iv_0_0_3,
       signal_data_iv_0_0_9,
       signal_data_iv_0_3_0,
       signal_data_iv_0_3_3,
       signal_data_iv_0_3_2,
       signal_data_iv_0_9_0,
       signal_data_iv_0_9_3,
       signal_data_iv_0_9_2,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_5,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_216,
       N_249,
       N_184,
       N_200,
       N_255,
       N_249_0,
       N_233,
       N_262,
       N_111,
       N_95,
       N_250,
       N_87,
       N_210,
       N_214,
       N_186,
       N_174,
       N_158,
       N_134,
       N_126,
       N_118,
       N_150,
       N_235,
       N_202,
       N_218,
       N_223
    );
output [14:14] addresult_RNI8MQ7;
input  [10:10] addresult_RNIFE5C;
input  [11:4] signal_data_0_iv_i_2;
input  [5:5] addresult_RNIBOIB;
output [11:4] signal_data_0_iv_i_5;
input  [1:1] signal_data_iv_0_0_3;
output [1:1] signal_data_iv_0_0_9;
input  signal_data_iv_0_3_0;
input  signal_data_iv_0_3_3;
input  signal_data_iv_0_3_2;
output signal_data_iv_0_9_0;
output signal_data_iv_0_9_3;
output signal_data_iv_0_9_2;
input  [4:0] un1_n_s_change_0_1;
input  [11:0] un1_ten_choice_one_0_5;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
output N_216;
input  N_249;
output N_184;
output N_200;
input  N_255;
input  N_249_0;
output N_233;
input  N_262;
output N_111;
output N_95;
input  N_250;
output N_87;
input  N_210;
input  N_214;
input  N_186;
input  N_174;
input  N_158;
input  N_134;
input  N_126;
input  N_118;
input  N_150;
input  N_235;
input  N_202;
input  N_218;
input  N_223;

    wire d_m5_0_0, d_N_8_0, d_m5_0_a4_0_0, \addresult_1[10] , 
        \addresult_1[9] , ADD_20x20_slow_I12_un1_CO1_m7, 
        ADD_20x20_slow_I12_un1_CO1_m1, ADD_20x20_slow_I12_un1_CO1_m7_2, 
        I8_un1_CO1, ADD_20x20_slow_I10_un1_CO1_0, 
        ADD_20x20_slow_I12_un1_CO1_m7_1, ADD_20x20_slow_I17_CO1_0, 
        \addresult_1[17] , ADD_20x20_slow_I16_un1_CO1_s, d_m6_i_0, 
        \addresult_1[11] , \addresult_1[12] , ADD_20x20_slow_I11_S_0_0, 
        d_m6_i_a4_0, ADD_20x20_slow_I8_S_0_0, \addresult_1[8] , 
        ADD_20x20_slow_I10_un1_CO1_0_m6_0, ADD_20x20_slow_I3_S_0_0, 
        \addresult_1[3] , d_m5_0_a4_0, 
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_1, 
        ADD_20x20_slow_I4_un1_CO1_0_N_12, ADD_20x20_slow_I2_un1_CO1_0, 
        N228, I2_un3_CO1_i, ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_1, 
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_0, \addresult_1[4] , 
        ADD_20x20_slow_I2_un3_CO1_m2_0_a2_0, \addresult_1[2] , 
        ADD_20x20_slow_I19_Y_0_m6_e_3, \addresult_1[13] , 
        ADD_20x20_slow_I19_Y_0_m6_e_0, ADD_20x20_slow_I19_Y_0_m6_e_2, 
        ADD_20x20_slow_I19_Y_0_m6_e_1, \addresult_1[15] , 
        \addresult_1[16] , \addresult_1[18] , \addresult_1[14] , N_217, 
        N_201, N_234, N_167, N_151, N_119, N_127, N_135, N_143, N_159, 
        N_175, N_185, N228_tz_tz, \addresult_RNIDQ8CC[10]_net_1 , 
        \addresult_RNIB4805[10]_net_1 , 
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_1, \addresult_1[1] , 
        \addresult_1[0] , \un3_addresult[10] , N244, 
        \un3_addresult[8] , N240, \un3_addresult[4] , N232, 
        \un3_addresult[3] , I2_un1_CO1, \un3_addresult[6] , 
        \addresult_1[6] , N236, \un3_addresult[1] , I0_un1_CO1, 
        \un3_addresult[2] , \un3_addresult[5] , \addresult_1[5] , 
        I4_un1_CO1, \un3_addresult[7] , \un1_add_reg_5_i[7] , 
        I6_un1_CO1_i, I2_un5_CO1_i, ADD_20x20_slow_I19_Y_0_m6_e_1_0, 
        ADD_20x20_slow_I10_un1_CO1_0_N_7_i, ADD_20x20_slow_I9_S_0_0, 
        \addresult_RNIKAD31[9]_net_1 , 
        ADD_20x20_slow_I4_un1_CO1_0_m8_i, 
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_o3_0, I14_un1_CO1, 
        I12_un1_CO1, \un3_addresult[11] , I10_un1_CO1, 
        \un3_addresult[9] , ADD_20x20_slow_I1_CO1_0_tz_tz_tz, 
        \addresult_RNIUG9P4[7]_net_1 , \addresult_RNO_1[19] , r_N_7_0, 
        \addresult_1[19] , \un3_addresult[12] , \un3_addresult[13] , 
        \un3_addresult[14] , \un3_addresult[18] , \un3_addresult[17] , 
        \un3_addresult[16] , \un3_addresult[15] , \un3_addresult[0] , 
        GND, VCC, GND_0, VCC_0;
    
    XOR2 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(I10_un1_CO1), .B(
        ADD_20x20_slow_I11_S_0_0), .Y(\un3_addresult[11] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[12] ));
    NOR3C \addresult_RNIU7L61[11]  (.A(N_151), .B(N_150), .C(
        signal_data_0_iv_i_2[11]), .Y(signal_data_0_iv_i_5[11]));
    OA1A \addresult_RNICIJ07[11]  (.A(\addresult_1[11] ), .B(
        un1_ten_choice_one_0_5[11]), .C(ADD_20x20_slow_I10_un1_CO1_0), 
        .Y(d_m6_i_a4_0));
    OR2 \addresult_RNI9MQ7[15]  (.A(\addresult_1[15] ), .B(N_250), .Y(
        N_111));
    XOR2 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        ADD_20x20_slow_I8_S_0_0), .B(N240), .Y(\un3_addresult[8] ));
    AO1C un3_addresult_ADD_20x20_slow_I1_CO1_tz_tz (.A(
        un1_n_s_change_0_1[1]), .B(ADD_20x20_slow_I1_CO1_0_tz_tz_tz), 
        .C(ADD_20x20_slow_I1_un5_CO1_m2_0_a2_1), .Y(N228_tz_tz));
    NOR3C \addresult_RNI8QUM1[1]  (.A(N_235), .B(N_234), .C(
        signal_data_iv_0_0_3[1]), .Y(signal_data_iv_0_0_9[1]));
    OR2 \addresult_RNI4MQ7[10]  (.A(\addresult_1[10] ), .B(N_250), .Y(
        N_143));
    NOR3C \addresult_RNIQ7L61[10]  (.A(N_143), .B(
        addresult_RNIFE5C[10]), .C(signal_data_0_iv_i_2[10]), .Y(
        signal_data_0_iv_i_5[10]));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[10] ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[6] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(I2_un1_CO1), .B(
        \addresult_1[3] ), .C(un1_ten_choice_one_0_5[3]), .Y(N232));
    OR2 \addresult_RNIMT97[9]  (.A(\addresult_1[9] ), .B(N_250), .Y(
        N_135));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[8] ));
    XOR2 un3_addresult_ADD_20x20_slow_I3_S_0_0 (.A(\addresult_1[3] ), 
        .B(un1_ten_choice_one_0_5[3]), .Y(ADD_20x20_slow_I3_S_0_0));
    OR2A \addresult_RNIVQCA_0[9]  (.A(un1_ten_choice_one_0_5[9]), .B(
        d_m5_0_a4_0_0), .Y(d_N_8_0));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un3_CO1_m2_0_a2_0 (.A(
        \addresult_1[2] ), .B(un1_n_s_change_0_1[2]), .Y(
        ADD_20x20_slow_I2_un3_CO1_m2_0_a2_0));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(I0_un1_CO1), .B(
        \addresult_1[1] ), .C(un1_ten_choice_one_0_5[1]), .Y(
        \un3_addresult[1] ));
    NOR3C \addresult_RNIM0JC1[5]  (.A(N_167), .B(addresult_RNIBOIB[5]), 
        .C(signal_data_0_iv_i_2[5]), .Y(signal_data_0_iv_i_5[5]));
    MX2C un3_addresult_ADD_20x20_slow_I10_un1_CO1_1 (.A(
        \addresult_RNIKAD31[9]_net_1 ), .B(
        \addresult_RNIUG9P4[7]_net_1 ), .S(
        ADD_20x20_slow_I10_un1_CO1_0_N_7_i), .Y(
        ADD_20x20_slow_I10_un1_CO1_0));
    AO1A un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_0_1 (.A(
        un1_n_s_change_0_1[3]), .B(\addresult_1[3] ), .C(
        \addresult_1[4] ), .Y(ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_0));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[15] ));
    XOR2 \addresult_RNO[19]  (.A(r_N_7_0), .B(\addresult_1[19] ), .Y(
        \addresult_RNO_1[19] ));
    OR2B un3_addresult_ADD_20x20_slow_I2_un1_CO1 (.A(
        ADD_20x20_slow_I2_un1_CO1_0), .B(I2_un5_CO1_i), .Y(I2_un1_CO1));
    VCC VCC_i (.Y(VCC));
    OR2B \addresult_RNI4FPB[3]  (.A(\addresult_1[3] ), .B(N_262), .Y(
        N_201));
    MAJ3 un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I4_un1_CO1), .B(
        \addresult_1[5] ), .C(un1_ten_choice_one_0_5[5]), .Y(N236));
    NOR3C un3_addresult_ADD_20x20_slow_I10_un1_CO1_0_m6 (.A(
        ADD_20x20_slow_I8_S_0_0), .B(ADD_20x20_slow_I10_un1_CO1_0_m6_0)
        , .C(ADD_20x20_slow_I9_S_0_0), .Y(
        ADD_20x20_slow_I10_un1_CO1_0_N_7_i));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_0 (.A(
        \addresult_1[18] ), .B(\addresult_1[14] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_0));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[4] ));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0_5[0]), .B(\addresult_1[0] ), .Y(
        \un3_addresult[0] ));
    OR2 \addresult_RNI7MQ7[13]  (.A(\addresult_1[13] ), .B(N_250), .Y(
        N_95));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[16] ));
    OR3A \addresult_RNIUVAC[16]  (.A(\addresult_1[16] ), .B(N_249), .C(
        N_255), .Y(N_184));
    NOR3C \addresult_RNI4IUM1[0]  (.A(N_186), .B(N_185), .C(
        signal_data_iv_0_3_0), .Y(signal_data_iv_0_9_0));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_5[5]), .B(\addresult_1[5] ), .C(
        I4_un1_CO1), .Y(\un3_addresult[5] ));
    MIN3 \addresult_RNIUG9P4[7]  (.A(I6_un1_CO1_i), .B(
        \un1_add_reg_5_i[7] ), .C(un1_ten_choice_one_0_5[7]), .Y(
        \addresult_RNIUG9P4[7]_net_1 ));
    OR2 \addresult_RNI6MQ7[12]  (.A(\addresult_1[12] ), .B(N_250), .Y(
        N_87));
    AX1C un3_addresult_ADD_20x20_slow_I14_S_0 (.A(I12_un1_CO1), .B(
        \addresult_1[13] ), .C(\addresult_1[14] ), .Y(
        \un3_addresult[14] ));
    XNOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0_5[4]), .B(\addresult_1[4] ), .C(N232), .Y(
        \un3_addresult[4] ));
    OR2A un3_addresult_ADD_20x20_slow_I2_un5_CO1 (.A(\addresult_1[2] ), 
        .B(N228), .Y(I2_un5_CO1_i));
    AX1C un3_addresult_ADD_20x20_slow_I18_S_0 (.A(I14_un1_CO1), .B(
        ADD_20x20_slow_I17_CO1_0), .C(\addresult_1[18] ), .Y(
        \un3_addresult[18] ));
    AO1A \addresult_RNIVQCA[9]  (.A(un1_ten_choice_one_0_5[9]), .B(
        \addresult_1[9] ), .C(\addresult_1[10] ), .Y(d_m5_0_a4_0));
    OAI1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i (.A(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_o3_0), .B(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_1), .C(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_1), .Y(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i));
    OR2 \addresult_RNI5MQ7[11]  (.A(\addresult_1[11] ), .B(N_250), .Y(
        N_151));
    AND2 \addresult_RNI5FLJ[9]  (.A(d_N_8_0), .B(
        un1_ten_choice_one_0_5[10]), .Y(d_m5_0_0));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[5] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_1[8] ), .C(un1_ten_choice_one_0_5[8]), .Y(
        I8_un1_CO1));
    NOR3C \addresult_RNIC2VM1[2]  (.A(N_218), .B(N_217), .C(
        signal_data_iv_0_3_2), .Y(signal_data_iv_0_9_2));
    AO13 \addresult_RNI0A6AC[11]  (.A(\addresult_1[11] ), .B(
        I10_un1_CO1), .C(un1_ten_choice_one_0_5[11]), .Y(r_N_7_0));
    OA1 un3_addresult_ADD_20x20_slow_I2_un1_CO1_0 (.A(N228), .B(
        un1_n_s_change_0_1[2]), .C(I2_un3_CO1_i), .Y(
        ADD_20x20_slow_I2_un1_CO1_0));
    OR2 \addresult_RNIID97[5]  (.A(\addresult_1[5] ), .B(N_250), .Y(
        N_167));
    OR2B \addresult_RNI13PB[0]  (.A(\addresult_1[0] ), .B(N_262), .Y(
        N_185));
    XNOR2 un3_addresult_ADD_20x20_slow_I12_un1_CO1_m1 (.A(
        un1_ten_choice_one_0_5[9]), .B(I8_un1_CO1), .Y(
        ADD_20x20_slow_I12_un1_CO1_m1));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[2] ));
    MIN3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1_i), .B(
        \un1_add_reg_5_i[7] ), .C(un1_ten_choice_one_0_5[7]), .Y(N240));
    NOR3C un3_addresult_ADD_20x20_slow_I14_un1_CO1 (.A(
        \addresult_1[13] ), .B(\addresult_1[14] ), .C(I12_un1_CO1), .Y(
        I14_un1_CO1));
    NOR3C \addresult_RNI61LC1[9]  (.A(N_135), .B(N_134), .C(
        signal_data_0_iv_i_2[9]), .Y(signal_data_0_iv_i_5[9]));
    OR2B \addresult_RNI3BPB[2]  (.A(\addresult_1[2] ), .B(N_262), .Y(
        N_217));
    OR3A \addresult_RNI10BC[19]  (.A(\addresult_1[19] ), .B(N_249_0), 
        .C(N_255), .Y(N_200));
    AO1A un3_addresult_ADD_20x20_slow_I1_CO1_0_tz_tz_tz (.A(
        un1_n_s_change_0_1[0]), .B(\addresult_1[0] ), .C(
        \addresult_1[1] ), .Y(ADD_20x20_slow_I1_CO1_0_tz_tz_tz));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e (.A(
        ADD_20x20_slow_I19_Y_0_m6_e_2), .B(
        ADD_20x20_slow_I19_Y_0_m6_e_1), .C(
        ADD_20x20_slow_I19_Y_0_m6_e_3), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_1_0));
    OR2 \addresult_RNILP97[8]  (.A(\addresult_1[8] ), .B(N_250), .Y(
        N_127));
    NOR3C \addresult_RNI2HKC1[8]  (.A(N_127), .B(N_126), .C(
        signal_data_0_iv_i_2[8]), .Y(signal_data_0_iv_i_5[8]));
    XOR2 un3_addresult_ADD_20x20_slow_I8_S_0_0 (.A(\addresult_1[8] ), 
        .B(un1_ten_choice_one_0_5[8]), .Y(ADD_20x20_slow_I8_S_0_0));
    AX1C un3_addresult_ADD_20x20_slow_I16_S_0 (.A(I14_un1_CO1), .B(
        \addresult_1[15] ), .C(\addresult_1[16] ), .Y(
        \un3_addresult[16] ));
    NOR2A un3_addresult_ADD_20x20_slow_I10_un1_CO1_0_m6_0 (.A(
        un1_ten_choice_one_0_5[10]), .B(\addresult_1[10] ), .Y(
        ADD_20x20_slow_I10_un1_CO1_0_m6_0));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[3] ));
    AND2 un3_addresult_ADD_20x20_slow_I12_un1_CO1_m7 (.A(
        ADD_20x20_slow_I12_un1_CO1_m1), .B(
        ADD_20x20_slow_I12_un1_CO1_m7_2), .Y(
        ADD_20x20_slow_I12_un1_CO1_m7));
    AX1C un3_addresult_ADD_20x20_slow_I17_S_0 (.A(
        ADD_20x20_slow_I16_un1_CO1_s), .B(I14_un1_CO1), .C(
        \addresult_1[17] ), .Y(\un3_addresult[17] ));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[14] ));
    OR3A un3_addresult_ADD_20x20_slow_I1_CO1 (.A(N228_tz_tz), .B(N_214)
        , .C(N_210), .Y(N228));
    XOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(r_N_7_0), .B(
        \addresult_1[12] ), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    AOI1B un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i_o3_0 (.A(
        un1_n_s_change_0_1[2]), .B(N228), .C(\addresult_1[2] ), .Y(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_o3_0));
    AO1B un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(\addresult_1[4] ), 
        .B(N232), .C(ADD_20x20_slow_I4_un1_CO1_0_m8_i), .Y(I4_un1_CO1));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_1 (.A(
        \addresult_1[15] ), .B(\addresult_1[16] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_1));
    OR2 \addresult_RNIJH97[6]  (.A(\addresult_1[6] ), .B(N_250), .Y(
        N_175));
    NOR3C \addresult_RNIIGIC1[4]  (.A(N_159), .B(N_158), .C(
        signal_data_0_iv_i_2[4]), .Y(signal_data_0_iv_i_5[4]));
    NOR3A un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i_1 (.A(
        ADD_20x20_slow_I4_un1_CO1_0_N_12), .B(un1_n_s_change_0_1[4]), 
        .C(N_223), .Y(ADD_20x20_slow_I4_un1_CO1_0_m8_i_1));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_2 (.A(
        \addresult_1[17] ), .B(\addresult_1[12] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_2));
    AND2 un3_addresult_ADD_20x20_slow_I12_un1_CO1_m7_2 (.A(
        ADD_20x20_slow_I10_un1_CO1_0), .B(
        ADD_20x20_slow_I12_un1_CO1_m7_1), .Y(
        ADD_20x20_slow_I12_un1_CO1_m7_2));
    XOR2 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(\addresult_1[15] ), 
        .B(I14_un1_CO1), .Y(\un3_addresult[15] ));
    OR2B \addresult_RNI27PB[1]  (.A(\addresult_1[1] ), .B(N_262), .Y(
        N_234));
    NOR3C un3_addresult_ADD_20x20_slow_I12_un1_CO1_m7_1 (.A(
        \addresult_1[10] ), .B(\addresult_1[12] ), .C(
        ADD_20x20_slow_I11_S_0_0), .Y(ADD_20x20_slow_I12_un1_CO1_m7_1));
    AO1B un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(
        \addresult_1[10] ), .B(N244), .C(ADD_20x20_slow_I10_un1_CO1_0), 
        .Y(I10_un1_CO1));
    AO1D un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_1 (.A(
        un1_n_s_change_0_1[2]), .B(N228), .C(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_0), .Y(
        ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_1));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[11] ));
    OR3B un3_addresult_ADD_20x20_slow_I1_un5_CO1_m2_0_a2_1 (.A(
        \addresult_1[1] ), .B(\addresult_1[0] ), .C(
        un1_n_s_change_0_1[0]), .Y(ADD_20x20_slow_I1_un5_CO1_m2_0_a2_1)
        );
    MX2A un3_addresult_ADD_20x20_slow_I12_un1_CO1_0 (.A(
        \addresult_RNIDQ8CC[10]_net_1 ), .B(\addresult_1[9] ), .S(
        ADD_20x20_slow_I12_un1_CO1_m7), .Y(I12_un1_CO1));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[17] ));
    AO13 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(\addresult_1[9] ), .B(
        I8_un1_CO1), .C(un1_ten_choice_one_0_5[9]), .Y(N244));
    NOR3C \addresult_RNIGAVM1[3]  (.A(N_202), .B(N_201), .C(
        signal_data_iv_0_3_3), .Y(signal_data_iv_0_9_3));
    OR3A \addresult_RNIVVAC[17]  (.A(\addresult_1[17] ), .B(N_249_0), 
        .C(N_255), .Y(N_233));
    OA1A \addresult_RNIM3DB[11]  (.A(un1_ten_choice_one_0_5[11]), .B(
        \addresult_1[11] ), .C(\addresult_1[12] ), .Y(d_m6_i_0));
    NOR2B un3_addresult_ADD_20x20_slow_I17_CO1_0 (.A(\addresult_1[17] )
        , .B(ADD_20x20_slow_I16_un1_CO1_s), .Y(
        ADD_20x20_slow_I17_CO1_0));
    OR3A \addresult_RNI00BC[18]  (.A(\addresult_1[18] ), .B(N_249), .C(
        N_255), .Y(N_216));
    OR3A un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_m8_i_a4_0 (.A(
        un1_n_s_change_0_1[3]), .B(\addresult_1[4] ), .C(
        \addresult_1[3] ), .Y(ADD_20x20_slow_I4_un1_CO1_0_N_12));
    AO1B \addresult_RNIDQ8CC[10]  (.A(d_m6_i_a4_0), .B(
        \addresult_RNIB4805[10]_net_1 ), .C(d_m6_i_0), .Y(
        \addresult_RNIDQ8CC[10]_net_1 ));
    MIN3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult_1[6] ), .C(un1_ten_choice_one_0_5[6]), .Y(
        I6_un1_CO1_i));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_5[10]), .B(\addresult_1[10] ), .C(N244), 
        .Y(\un3_addresult[10] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I9_S_0_0 (.A(
        un1_ten_choice_one_0_5[9]), .B(\addresult_1[9] ), .Y(
        ADD_20x20_slow_I9_S_0_0));
    DFN1P0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        \un1_add_reg_5_i[7] ));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_3 (.A(
        \addresult_1[13] ), .B(ADD_20x20_slow_I19_Y_0_m6_e_0), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_3));
    OR2A \addresult_RNIKL97[7]  (.A(\un1_add_reg_5_i[7] ), .B(N_250), 
        .Y(N_119));
    OA1 \addresult_RNIKAD31[9]  (.A(un1_ten_choice_one_0_5[8]), .B(
        d_m5_0_a4_0), .C(d_m5_0_0), .Y(\addresult_RNIKAD31[9]_net_1 ));
    XOR2 un3_addresult_ADD_20x20_slow_I13_S_0 (.A(\addresult_1[13] ), 
        .B(I12_un1_CO1), .Y(\un3_addresult[13] ));
    OR2 \addresult_RNIUMJ1[9]  (.A(\addresult_1[10] ), .B(
        \addresult_1[9] ), .Y(d_m5_0_a4_0_0));
    XOR2 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        ADD_20x20_slow_I3_S_0_0), .B(I2_un1_CO1), .Y(
        \un3_addresult[3] ));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[18] ));
    NOR2B un3_addresult_ADD_20x20_slow_I16_un1_CO1_s (.A(
        \addresult_1[16] ), .B(\addresult_1[15] ), .Y(
        ADD_20x20_slow_I16_un1_CO1_s));
    XOR3 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        un1_ten_choice_one_0_5[6]), .B(\addresult_1[6] ), .C(N236), .Y(
        \un3_addresult[6] ));
    OR2B \addresult_RNIB4805[10]  (.A(\addresult_1[10] ), .B(
        I8_un1_CO1), .Y(\addresult_RNIB4805[10]_net_1 ));
    NOR3C \addresult_RNIQGJC1[6]  (.A(N_175), .B(N_174), .C(
        signal_data_0_iv_i_2[6]), .Y(signal_data_0_iv_i_5[6]));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[13] ));
    NOR3C \addresult_RNIU0KC1[7]  (.A(N_119), .B(N_118), .C(
        signal_data_0_iv_i_2[7]), .Y(signal_data_0_iv_i_5[7]));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[9] ));
    DFN1E1C0 \addresult[19]  (.D(\addresult_RNO_1[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .E(
        ADD_20x20_slow_I19_Y_0_m6_e_1_0), .Q(\addresult_1[19] ));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[0] ));
    OR2B un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(
        un1_ten_choice_one_0_5[0]), .B(\addresult_1[0] ), .Y(
        I0_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0_5[7]), .B(\un1_add_reg_5_i[7] ), .C(
        I6_un1_CO1_i), .Y(\un3_addresult[7] ));
    XOR2 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(I8_un1_CO1), .B(
        ADD_20x20_slow_I9_S_0_0), .Y(\un3_addresult[9] ));
    XOR3 un3_addresult_ADD_20x20_slow_I2_S_0 (.A(N228), .B(
        \addresult_1[2] ), .C(un1_ten_choice_one_0_5[2]), .Y(
        \un3_addresult[2] ));
    OR2 \addresult_RNIH997[4]  (.A(\addresult_1[4] ), .B(N_250), .Y(
        N_159));
    VCC VCC_i_0 (.Y(VCC_0));
    OR3A un3_addresult_ADD_20x20_slow_I2_un3_CO1_m2_0_a2 (.A(
        ADD_20x20_slow_I2_un3_CO1_m2_0_a2_0), .B(N_214), .C(N_210), .Y(
        I2_un3_CO1_i));
    XNOR2 un3_addresult_ADD_20x20_slow_I11_S_0_0 (.A(
        un1_ten_choice_one_0_5[11]), .B(\addresult_1[11] ), .Y(
        ADD_20x20_slow_I11_S_0_0));
    GND GND_i_0 (.Y(GND_0));
    OR2 \addresult_RNI8MQ7[14]  (.A(\addresult_1[14] ), .B(N_250), .Y(
        addresult_RNI8MQ7[14]));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[1] ));
    
endmodule


module add_reg_add_reg_2_4(
       un1_n_s_change_0_1,
       signal_data_0_iv_i_5,
       signal_data_0_iv_i_3,
       signal_data_0_iv_i_0,
       signal_data_iv_0_0_10,
       signal_data_iv_0_0_6,
       signal_data_iv_0_0_13,
       signal_data_iv_0_10_0,
       signal_data_iv_0_10_3,
       signal_data_iv_0_10_2,
       signal_data_iv_0_6_0,
       signal_data_iv_0_6_3,
       signal_data_iv_0_6_2,
       signal_data_iv_0_13_0,
       signal_data_iv_0_13_3,
       signal_data_iv_0_13_2,
       un1_ten_choice_one_0,
       addresult_4_10,
       addresult_4_8,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_226,
       N_249,
       N_194,
       N_210,
       N_254,
       N_249_0,
       N_243,
       N_108,
       N_92,
       N_222,
       N_25_i_0,
       N_20_i_0,
       N_12_i_0,
       N_14_i_0,
       N_16_i_0,
       N_18_i_0,
       N_22_i_0,
       N_27_i_0,
       N_196,
       N_39,
       N_245,
       N_212,
       N_228,
       N_271
    );
input  [2:0] un1_n_s_change_0_1;
input  [11:4] signal_data_0_iv_i_5;
input  [11:4] signal_data_0_iv_i_3;
input  [11:4] signal_data_0_iv_i_0;
input  [1:1] signal_data_iv_0_0_10;
input  [1:1] signal_data_iv_0_0_6;
output [1:1] signal_data_iv_0_0_13;
input  signal_data_iv_0_10_0;
input  signal_data_iv_0_10_3;
input  signal_data_iv_0_10_2;
input  signal_data_iv_0_6_0;
input  signal_data_iv_0_6_3;
input  signal_data_iv_0_6_2;
output signal_data_iv_0_13_0;
output signal_data_iv_0_13_3;
output signal_data_iv_0_13_2;
input  [11:0] un1_ten_choice_one_0;
output addresult_4_10;
output addresult_4_8;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
output N_226;
input  N_249;
output N_194;
output N_210;
input  N_254;
input  N_249_0;
output N_243;
output N_108;
output N_92;
input  N_222;
output N_25_i_0;
output N_20_i_0;
output N_12_i_0;
output N_14_i_0;
output N_16_i_0;
output N_18_i_0;
output N_22_i_0;
output N_27_i_0;
input  N_196;
input  N_39;
input  N_245;
input  N_212;
input  N_228;
input  N_271;

    wire ADD_20x20_slow_I18_un1_CO1_1, \addresult_5[17] , 
        \addresult_5[18] , \addresult_5[16] , ADD_20x20_slow_I17_CO1_0, 
        ADD_20x20_slow_I5_CO1_0_tz_0, \addresult_5[4] , N232, 
        \addresult_4[5] , d_m5_i_0, \addresult_5[14] , 
        \addresult_5[12] , ADD_20x20_slow_I14_un1_CO1_m6_1, 
        \addresult_5[10] , \signal_data_iv_0_7[2] , \addresult_5[2] , 
        \signal_data_iv_0_7[3] , \addresult_5[3] , 
        \signal_data_iv_0_0_7[1] , \addresult_5[1] , 
        \signal_data_0_iv_i_4[5] , \signal_data_0_iv_i_4[11] , 
        \addresult_5[11] , \signal_data_0_iv_i_4[7] , \addresult_4[7] , 
        \signal_data_0_iv_i_4[8] , \addresult_5[8] , 
        \signal_data_0_iv_i_4[9] , \un1_add_reg_0_i[9] , 
        \signal_data_0_iv_i_4[10] , \signal_data_0_iv_i_4[4] , 
        \signal_data_0_iv_i_4[6] , \addresult_5[6] , 
        \signal_data_iv_0_7[0] , \addresult_5[0] , 
        \addresult_RNIQ2OC1[11]_net_1 , d_N_8_1, d_N_7_1, 
        ADD_20x20_slow_I14_un1_CO1_N_7_i, \un3_addresult[10] , N244, 
        \un3_addresult[9] , I8_un1_CO1_i, \un3_addresult[8] , N240, 
        \un3_addresult[7] , I6_un1_CO1, \un3_addresult[6] , N236, 
        \un3_addresult[5] , I4_un1_CO1, \un3_addresult[4] , 
        \un3_addresult[3] , I2_un1_CO1, \un3_addresult[2] , N228, 
        \un3_addresult[1] , I0_un1_CO1, \un3_addresult[11] , 
        I10_un1_CO1, ADD_20x20_slow_I1_CO1_0_tz, I14_un1_CO1, 
        \addresult_RNIFBP77[9]_net_1 , I1_un3_CO1, 
        ADD_20x20_slow_I2_un1_CO1_N_7, ADD_20x20_slow_I2_un1_CO1_N_4, 
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_0, ADD_20x20_slow_I5_CO1_0, 
        ADD_20x20_slow_I4_un1_CO1_0, I5_un5_CO1, N248, I12_un1_CO1, 
        N262, \un3_addresult[12] , \un3_addresult[13] , 
        \un3_addresult[14] , \un3_addresult[15] , \un3_addresult[16] , 
        \un3_addresult[17] , \un3_addresult[18] , \un3_addresult[19] , 
        \addresult_5[19] , \un3_addresult[0] , GND, VCC, GND_0, VCC_0;
    
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(\addresult_5[11] ), 
        .B(un1_ten_choice_one_0[11]), .C(I10_un1_CO1), .Y(
        \un3_addresult[11] ));
    OR3A \addresult_RNIA6LE[19]  (.A(\addresult_5[19] ), .B(N_249_0), 
        .C(N_254), .Y(N_210));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[12] ));
    AOI1B \addresult_RNIU9BR[3]  (.A(\addresult_5[3] ), .B(N_271), .C(
        N_212), .Y(\signal_data_iv_0_7[3] ));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0[8]), .B(\addresult_5[8] ), .C(N240), .Y(
        \un3_addresult[8] ));
    OR2 \addresult_RNIFS4A[12]  (.A(\addresult_5[12] ), .B(N_39), .Y(
        N_92));
    NOR3C \addresult_RNIOLFR2[9]  (.A(\signal_data_0_iv_i_4[9] ), .B(
        signal_data_0_iv_i_3[9]), .C(signal_data_0_iv_i_5[9]), .Y(
        N_16_i_0));
    NOR3C \addresult_RNIG1214[0]  (.A(\signal_data_iv_0_7[0] ), .B(
        signal_data_iv_0_6_0), .C(signal_data_iv_0_10_0), .Y(
        signal_data_iv_0_13_0));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[10] ));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m7 (.A(N_222), .B(
        ADD_20x20_slow_I2_un1_CO1_N_7), .Y(I2_un1_CO1));
    NOR3C \addresult_RNIOKBR2[5]  (.A(\signal_data_0_iv_i_4[5] ), .B(
        signal_data_0_iv_i_3[5]), .C(signal_data_0_iv_i_5[5]), .Y(
        N_25_i_0));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[6] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(I2_un1_CO1), .B(
        \addresult_5[3] ), .C(un1_ten_choice_one_0[3]), .Y(N232));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[8] ));
    OR2 \addresult_RNIHS4A[14]  (.A(\addresult_5[14] ), .B(N_39), .Y(
        N_108));
    NOR3C \addresult_RNI0LCR2[6]  (.A(\signal_data_0_iv_i_4[6] ), .B(
        signal_data_0_iv_i_3[6]), .C(signal_data_0_iv_i_5[6]), .Y(
        N_27_i_0));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(
        un1_ten_choice_one_0[1]), .B(\addresult_5[1] ), .C(I0_un1_CO1), 
        .Y(\un3_addresult[1] ));
    OR2A un3_addresult_ADD_20x20_slow_I1_un3_CO1 (.A(I0_un1_CO1), .B(
        un1_n_s_change_0_1[1]), .Y(I1_un3_CO1));
    NOR3C \addresult_RNI02314[2]  (.A(\signal_data_iv_0_7[2] ), .B(
        signal_data_iv_0_6_2), .C(signal_data_iv_0_10_2), .Y(
        signal_data_iv_0_13_2));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_4_10));
    VCC VCC_i (.Y(VCC));
    AO1B un3_addresult_ADD_20x20_slow_I5_CO1_0 (.A(
        ADD_20x20_slow_I5_CO1_0_tz_0), .B(ADD_20x20_slow_I4_un1_CO1_0), 
        .C(un1_ten_choice_one_0[5]), .Y(ADD_20x20_slow_I5_CO1_0));
    OR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1tt_m1_e (.A(
        \addresult_5[0] ), .B(un1_n_s_change_0_1[0]), .Y(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_0));
    MAJ3 un3_addresult_ADD_20x20_slow_I11_CO1 (.A(I10_un1_CO1), .B(
        \addresult_5[11] ), .C(un1_ten_choice_one_0[11]), .Y(N248));
    OR2B un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I5_un5_CO1), .B(
        ADD_20x20_slow_I5_CO1_0), .Y(N236));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[4] ));
    NOR2A un3_addresult_ADD_20x20_slow_I15_CO1 (.A(addresult_4_10), .B(
        I14_un1_CO1), .Y(N262));
    NOR2B un3_addresult_ADD_20x20_slow_I12_un1_CO1 (.A(
        \addresult_5[12] ), .B(N248), .Y(I12_un1_CO1));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0[0]), .B(\addresult_5[0] ), .Y(
        \un3_addresult[0] ));
    AO18 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m6 (.A(
        ADD_20x20_slow_I2_un1_CO1_N_4), .B(un1_n_s_change_0_1[2]), .C(
        \addresult_5[2] ), .Y(ADD_20x20_slow_I2_un1_CO1_N_7));
    OR3A \addresult_RNI76LE[16]  (.A(\addresult_5[16] ), .B(N_249), .C(
        N_254), .Y(N_194));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[16] ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0[5]), .B(\addresult_4[5] ), .C(I4_un1_CO1), 
        .Y(\un3_addresult[5] ));
    AO1 \addresult_RNIDMTL[11]  (.A(un1_ten_choice_one_0[11]), .B(
        \addresult_5[11] ), .C(un1_ten_choice_one_0[10]), .Y(d_N_7_1));
    NOR3C \addresult_RNI8I314[3]  (.A(\signal_data_iv_0_7[3] ), .B(
        signal_data_iv_0_6_3), .C(signal_data_iv_0_10_3), .Y(
        signal_data_iv_0_13_3));
    AX1C un3_addresult_ADD_20x20_slow_I14_S_0 (.A(I12_un1_CO1), .B(
        addresult_4_8), .C(\addresult_5[14] ), .Y(\un3_addresult[14] ));
    NOR3C \addresult_RNIGM4N2[10]  (.A(\signal_data_0_iv_i_4[10] ), .B(
        signal_data_0_iv_i_3[10]), .C(signal_data_0_iv_i_5[10]), .Y(
        N_18_i_0));
    XOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0[4]), .B(\addresult_5[4] ), .C(N232), .Y(
        \un3_addresult[4] ));
    AX1C un3_addresult_ADD_20x20_slow_I18_S_0 (.A(N262), .B(
        ADD_20x20_slow_I17_CO1_0), .C(\addresult_5[18] ), .Y(
        \un3_addresult[18] ));
    OR3A \addresult_RNI86LE[17]  (.A(\addresult_5[17] ), .B(N_249_0), 
        .C(N_254), .Y(N_243));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[5] ));
    MIN3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_5[8] ), .C(un1_ten_choice_one_0[8]), .Y(
        I8_un1_CO1_i));
    AX1C un3_addresult_ADD_20x20_slow_I19_Y_0 (.A(N262), .B(
        ADD_20x20_slow_I18_un1_CO1_1), .C(\addresult_5[19] ), .Y(
        \un3_addresult[19] ));
    OA1 \addresult_RNIJS7M[8]  (.A(N_39), .B(\addresult_5[8] ), .C(
        signal_data_0_iv_i_0[8]), .Y(\signal_data_0_iv_i_4[8] ));
    OR2 \addresult_RNI72LC[11]  (.A(un1_ten_choice_one_0[11]), .B(
        \addresult_5[11] ), .Y(d_N_8_1));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[2] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult_4[7] ), .C(un1_ten_choice_one_0[7]), .Y(N240));
    AO18 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m3 (.A(
        un1_n_s_change_0_1[1]), .B(\addresult_5[1] ), .C(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_0), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_4));
    OR2B un3_addresult_ADD_20x20_slow_I5_un5_CO1 (.A(\addresult_4[5] ), 
        .B(I4_un1_CO1), .Y(I5_un5_CO1));
    NOR3C \addresult_RNIQ2OC1[11]  (.A(d_N_8_1), .B(d_m5_i_0), .C(
        d_N_7_1), .Y(\addresult_RNIQ2OC1[11]_net_1 ));
    XOR2 un3_addresult_ADD_20x20_slow_I16_S_0 (.A(\addresult_5[16] ), 
        .B(N262), .Y(\un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[3] ));
    AOI1B \addresult_RNIOTAR[0]  (.A(\addresult_5[0] ), .B(N_271), .C(
        N_196), .Y(\signal_data_iv_0_7[0] ));
    XA1 un3_addresult_ADD_20x20_slow_I14_un1_CO1_m6 (.A(
        \addresult_5[11] ), .B(un1_ten_choice_one_0[11]), .C(
        ADD_20x20_slow_I14_un1_CO1_m6_1), .Y(
        ADD_20x20_slow_I14_un1_CO1_N_7_i));
    AX1C un3_addresult_ADD_20x20_slow_I17_S_0 (.A(N262), .B(
        \addresult_5[16] ), .C(\addresult_5[17] ), .Y(
        \un3_addresult[17] ));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[14] ));
    AO1B un3_addresult_ADD_20x20_slow_I1_CO1 (.A(\addresult_5[1] ), .B(
        ADD_20x20_slow_I1_CO1_0_tz), .C(I1_un3_CO1), .Y(N228));
    XOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(\addresult_5[12] ), 
        .B(N248), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    NOR3C \addresult_RNIOH214[1]  (.A(\signal_data_iv_0_0_7[1] ), .B(
        signal_data_iv_0_0_6[1]), .C(signal_data_iv_0_0_10[1]), .Y(
        signal_data_iv_0_0_13[1]));
    AO1B un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(\addresult_5[4] ), 
        .B(N232), .C(ADD_20x20_slow_I4_un1_CO1_0), .Y(I4_un1_CO1));
    NOR3C \addresult_RNIGLER2[8]  (.A(\signal_data_0_iv_i_4[8] ), .B(
        signal_data_0_iv_i_3[8]), .C(signal_data_0_iv_i_5[8]), .Y(
        N_14_i_0));
    OA1 \addresult_RNIRC5N[10]  (.A(N_39), .B(\addresult_5[10] ), .C(
        signal_data_0_iv_i_0[10]), .Y(\signal_data_0_iv_i_4[10] ));
    OR3A \addresult_RNI96LE[18]  (.A(\addresult_5[18] ), .B(N_249), .C(
        N_254), .Y(N_226));
    OA1 \addresult_RNITC5N[11]  (.A(N_39), .B(\addresult_5[11] ), .C(
        signal_data_0_iv_i_0[11]), .Y(\signal_data_0_iv_i_4[11] ));
    OA1A \addresult_RNIL48M[9]  (.A(\un1_add_reg_0_i[9] ), .B(N_39), 
        .C(signal_data_0_iv_i_0[9]), .Y(\signal_data_0_iv_i_4[9] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(addresult_4_10), .B(
        I14_un1_CO1), .Y(\un3_addresult[15] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult_5[10] ), .C(un1_ten_choice_one_0[10]), .Y(
        I10_un1_CO1));
    AOI1B \addresult_RNIS5BR[2]  (.A(\addresult_5[2] ), .B(N_271), .C(
        N_228), .Y(\signal_data_iv_0_7[2] ));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[11] ));
    XA1 un3_addresult_ADD_20x20_slow_I14_un1_CO1_m6_1 (.A(
        un1_ten_choice_one_0[10]), .B(\addresult_5[10] ), .C(d_m5_i_0), 
        .Y(ADD_20x20_slow_I14_un1_CO1_m6_1));
    OA1 \addresult_RNID47M[5]  (.A(N_39), .B(\addresult_4[5] ), .C(
        signal_data_0_iv_i_0[5]), .Y(\signal_data_0_iv_i_4[5] ));
    OAI1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0 (.A(N232), .B(
        \addresult_5[4] ), .C(un1_ten_choice_one_0[4]), .Y(
        ADD_20x20_slow_I4_un1_CO1_0));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[17] ));
    MIN3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1_i), .B(
        \un1_add_reg_0_i[9] ), .C(un1_ten_choice_one_0[9]), .Y(N244));
    MIN3 \addresult_RNIFBP77[9]  (.A(I8_un1_CO1_i), .B(
        \un1_add_reg_0_i[9] ), .C(un1_ten_choice_one_0[9]), .Y(
        \addresult_RNIFBP77[9]_net_1 ));
    AOI1 un3_addresult_ADD_20x20_slow_I5_CO1_0_tz_0 (.A(
        \addresult_5[4] ), .B(N232), .C(\addresult_4[5] ), .Y(
        ADD_20x20_slow_I5_CO1_0_tz_0));
    NOR3C \addresult_RNIGKAR2[4]  (.A(\signal_data_0_iv_i_4[4] ), .B(
        signal_data_0_iv_i_3[4]), .C(signal_data_0_iv_i_5[4]), .Y(
        N_22_i_0));
    NOR2B un3_addresult_ADD_20x20_slow_I17_CO1_0 (.A(\addresult_5[17] )
        , .B(\addresult_5[16] ), .Y(ADD_20x20_slow_I17_CO1_0));
    OR2 un3_addresult_ADD_20x20_slow_I1_CO1_0_tz (.A(
        un1_ten_choice_one_0[1]), .B(I0_un1_CO1), .Y(
        ADD_20x20_slow_I1_CO1_0_tz));
    AOI1B \addresult_RNIQ1BR[1]  (.A(\addresult_5[1] ), .B(N_271), .C(
        N_245), .Y(\signal_data_iv_0_0_7[1] ));
    NOR3C \addresult_RNI6A5A[14]  (.A(addresult_4_8), .B(
        \addresult_5[14] ), .C(\addresult_5[12] ), .Y(d_m5_i_0));
    MAJ3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult_5[6] ), .C(un1_ten_choice_one_0[6]), .Y(I6_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0[10]), .B(\addresult_5[10] ), .C(N244), .Y(
        \un3_addresult[10] ));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[7] ));
    XOR2 un3_addresult_ADD_20x20_slow_I13_S_0 (.A(addresult_4_8), .B(
        I12_un1_CO1), .Y(\un3_addresult[13] ));
    XOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        un1_ten_choice_one_0[3]), .B(\addresult_5[3] ), .C(I2_un1_CO1), 
        .Y(\un3_addresult[3] ));
    OA1 \addresult_RNIFC7M[6]  (.A(N_39), .B(\addresult_5[6] ), .C(
        signal_data_0_iv_i_0[6]), .Y(\signal_data_0_iv_i_4[6] ));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[18] ));
    OA1 \addresult_RNIHK7M[7]  (.A(N_39), .B(\addresult_4[7] ), .C(
        signal_data_0_iv_i_0[7]), .Y(\signal_data_0_iv_i_4[7] ));
    XOR3 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        un1_ten_choice_one_0[6]), .B(\addresult_5[6] ), .C(N236), .Y(
        \un3_addresult[6] ));
    OA1 \addresult_RNIBS6M[4]  (.A(N_39), .B(\addresult_5[4] ), .C(
        signal_data_0_iv_i_0[4]), .Y(\signal_data_0_iv_i_4[4] ));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_4_8));
    NOR3C un3_addresult_ADD_20x20_slow_I18_un1_CO1_1 (.A(
        \addresult_5[17] ), .B(\addresult_5[18] ), .C(
        \addresult_5[16] ), .Y(ADD_20x20_slow_I18_un1_CO1_1));
    NOR3C \addresult_RNIOM4N2[11]  (.A(\signal_data_0_iv_i_4[11] ), .B(
        signal_data_0_iv_i_3[11]), .C(signal_data_0_iv_i_5[11]), .Y(
        N_20_i_0));
    MX2C un3_addresult_ADD_20x20_slow_I14_un1_CO1_0 (.A(
        \addresult_RNIQ2OC1[11]_net_1 ), .B(
        \addresult_RNIFBP77[9]_net_1 ), .S(
        ADD_20x20_slow_I14_un1_CO1_N_7_i), .Y(I14_un1_CO1));
    NOR3C \addresult_RNI8LDR2[7]  (.A(\signal_data_0_iv_i_4[7] ), .B(
        signal_data_0_iv_i_3[7]), .C(signal_data_0_iv_i_5[7]), .Y(
        N_12_i_0));
    DFN1P0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        \un1_add_reg_0_i[9] ));
    DFN1C0 \addresult[19]  (.D(\un3_addresult[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[19] ));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[0] ));
    NOR2B un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(
        un1_ten_choice_one_0[0]), .B(\addresult_5[0] ), .Y(I0_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0[7]), .B(\addresult_4[7] ), .C(I6_un1_CO1), 
        .Y(\un3_addresult[7] ));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0[9]), .B(\un1_add_reg_0_i[9] ), .C(
        I8_un1_CO1_i), .Y(\un3_addresult[9] ));
    XNOR3 un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        un1_ten_choice_one_0[2]), .B(\addresult_5[2] ), .C(N228), .Y(
        \un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[1] ));
    
endmodule


module ten_choice_one(
       un1_ten_choice_one_0_7_0,
       un1_ten_choice_one_0_7_2,
       un1_ten_choice_one_0_7_11,
       un1_ten_choice_one_0_7_10,
       un1_ten_choice_one_0_7_9,
       un1_ten_choice_one_0_7_8,
       un1_ten_choice_one_0_7_7,
       un1_ten_choice_one_0_7_6,
       un1_ten_choice_one_0_7_5,
       un1_ten_choice_one_0_7_3,
       un1_ten_choice_one_0_4_3,
       un1_ten_choice_one_0_4_1,
       un1_ten_choice_one_0_4_0,
       un1_ten_choice_one_0_4_11,
       un1_ten_choice_one_0_4_10,
       un1_ten_choice_one_0_4_9,
       un1_ten_choice_one_0_4_8,
       un1_ten_choice_one_0_4_7,
       un1_ten_choice_one_0_4_6,
       un1_ten_choice_one_0_4_5,
       un1_ten_choice_one_0_4_4,
       un1_ten_choice_one_0_3_1,
       un1_ten_choice_one_0_3_0,
       un1_ten_choice_one_0_3_10,
       un1_ten_choice_one_0_3_11,
       un1_ten_choice_one_0_3_9,
       un1_ten_choice_one_0_3_8,
       un1_ten_choice_one_0_3_7,
       un1_ten_choice_one_0_3_6,
       un1_ten_choice_one_0_3_5,
       un1_ten_choice_one_0_3_4,
       un1_ten_choice_one_0_3_3,
       un1_ten_choice_one_0,
       un1_ten_choice_one_0_6,
       un1_ten_choice_one_0_5,
       un1_ten_choice_one_0_1_2,
       un1_ten_choice_one_0_1_1,
       un1_ten_choice_one_0_1_0,
       un1_ten_choice_one_0_1_8,
       un1_ten_choice_one_0_1_10,
       un1_ten_choice_one_0_1_11,
       un1_ten_choice_one_0_1_9,
       un1_ten_choice_one_0_1_7,
       un1_ten_choice_one_0_1_6,
       un1_ten_choice_one_0_1_5,
       un1_ten_choice_one_0_1_4,
       addrout,
       dataeight_0_a2_0_0,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_2_0,
       un1_ten_choice_one_0_2_10,
       un1_ten_choice_one_0_2_9,
       un1_ten_choice_one_0_2_8,
       un1_ten_choice_one_0_2_7,
       un1_ten_choice_one_0_2_6,
       un1_ten_choice_one_0_2_5,
       un1_ten_choice_one_0_2_4,
       un1_ten_choice_one_0_2_3,
       un1_ten_choice_one_0_2_2,
       N_214,
       N_212,
       N_211,
       N_217,
       N_219,
       N_222,
       N_221,
       N_223,
       N_224,
       N_216,
       N_213,
       N_220,
       N_210,
       N_215
    );
output un1_ten_choice_one_0_7_0;
output un1_ten_choice_one_0_7_2;
output un1_ten_choice_one_0_7_11;
output un1_ten_choice_one_0_7_10;
output un1_ten_choice_one_0_7_9;
output un1_ten_choice_one_0_7_8;
output un1_ten_choice_one_0_7_7;
output un1_ten_choice_one_0_7_6;
output un1_ten_choice_one_0_7_5;
output un1_ten_choice_one_0_7_3;
output un1_ten_choice_one_0_4_3;
output un1_ten_choice_one_0_4_1;
output un1_ten_choice_one_0_4_0;
output un1_ten_choice_one_0_4_11;
output un1_ten_choice_one_0_4_10;
output un1_ten_choice_one_0_4_9;
output un1_ten_choice_one_0_4_8;
output un1_ten_choice_one_0_4_7;
output un1_ten_choice_one_0_4_6;
output un1_ten_choice_one_0_4_5;
output un1_ten_choice_one_0_4_4;
output un1_ten_choice_one_0_3_1;
output un1_ten_choice_one_0_3_0;
output un1_ten_choice_one_0_3_10;
output un1_ten_choice_one_0_3_11;
output un1_ten_choice_one_0_3_9;
output un1_ten_choice_one_0_3_8;
output un1_ten_choice_one_0_3_7;
output un1_ten_choice_one_0_3_6;
output un1_ten_choice_one_0_3_5;
output un1_ten_choice_one_0_3_4;
output un1_ten_choice_one_0_3_3;
output [11:0] un1_ten_choice_one_0;
output [11:1] un1_ten_choice_one_0_6;
output [11:0] un1_ten_choice_one_0_5;
output un1_ten_choice_one_0_1_2;
output un1_ten_choice_one_0_1_1;
output un1_ten_choice_one_0_1_0;
output un1_ten_choice_one_0_1_8;
output un1_ten_choice_one_0_1_10;
output un1_ten_choice_one_0_1_11;
output un1_ten_choice_one_0_1_9;
output un1_ten_choice_one_0_1_7;
output un1_ten_choice_one_0_1_6;
output un1_ten_choice_one_0_1_5;
output un1_ten_choice_one_0_1_4;
input  [3:0] addrout;
output [0:0] dataeight_0_a2_0_0;
input  [11:0] un1_n_s_change_0_1;
output un1_ten_choice_one_0_2_0;
output un1_ten_choice_one_0_2_10;
output un1_ten_choice_one_0_2_9;
output un1_ten_choice_one_0_2_8;
output un1_ten_choice_one_0_2_7;
output un1_ten_choice_one_0_2_6;
output un1_ten_choice_one_0_2_5;
output un1_ten_choice_one_0_2_4;
output un1_ten_choice_one_0_2_3;
output un1_ten_choice_one_0_2_2;
output N_214;
output N_212;
output N_211;
output N_217;
output N_219;
output N_222;
output N_221;
output N_223;
output N_224;
output N_216;
output N_213;
output N_220;
output N_210;
output N_215;

    wire GND, VCC, GND_0, VCC_0;
    
    OR2 \datasix_0_a2[1]  (.A(un1_n_s_change_0_1[1]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[1]));
    OR2 \datasix_0_a2_0[0]  (.A(N_214), .B(N_210), .Y(N_223));
    NOR2A \dataone_0_a2[3]  (.A(N_222), .B(un1_n_s_change_0_1[3]), .Y(
        un1_ten_choice_one_0[3]));
    NOR2A \datafive_0_a2[10]  (.A(N_217), .B(un1_n_s_change_0_1[10]), 
        .Y(un1_ten_choice_one_0_4_10));
    OR2 \dataeight_0_a2[2]  (.A(un1_n_s_change_0_1[2]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_2));
    NOR2 \datasix_0_a2[3]  (.A(un1_n_s_change_0_1[3]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[3]));
    OR2 \dataseven_0_a2[1]  (.A(un1_n_s_change_0_1[1]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[1]));
    NOR2A \datafive_0_a2[8]  (.A(N_217), .B(un1_n_s_change_0_1[8]), .Y(
        un1_ten_choice_one_0_4_8));
    NOR2A \datatwo_0_a2[10]  (.A(N_216), .B(un1_n_s_change_0_1[10]), 
        .Y(un1_ten_choice_one_0_1_10));
    OR2 \datasix_0_a2[4]  (.A(un1_n_s_change_0_1[4]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[4]));
    OR2 \dataseven_0_a2_0[0]  (.A(N_212), .B(N_210), .Y(N_221));
    NOR2 \dataseven_0_a2[11]  (.A(un1_n_s_change_0_1[11]), .B(N_221), 
        .Y(un1_ten_choice_one_0_6[11]));
    OR2A \datafive_0_a2[3]  (.A(N_217), .B(un1_n_s_change_0_1[3]), .Y(
        un1_ten_choice_one_0_4_3));
    OR2 \datatwo_0_a2_2[0]  (.A(addrout[2]), .B(addrout[0]), .Y(N_213));
    NOR2A \datatwo_0_a2[9]  (.A(N_216), .B(un1_n_s_change_0_1[9]), .Y(
        un1_ten_choice_one_0_1_9));
    NOR2 \dataseven_0_a2[3]  (.A(un1_n_s_change_0_1[3]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[3]));
    NOR2A \dataone_0_a2[0]  (.A(N_222), .B(un1_n_s_change_0_1[0]), .Y(
        un1_ten_choice_one_0[0]));
    OR2 \dataseven_0_a2[2]  (.A(un1_n_s_change_0_1[2]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[2]));
    NOR2A \datathree_0_a2[8]  (.A(N_224), .B(un1_n_s_change_0_1[8]), 
        .Y(un1_ten_choice_one_0_2_7));
    OR2 \datasix_0_a2[2]  (.A(un1_n_s_change_0_1[2]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[2]));
    NOR2A \datatwo_0_a2[7]  (.A(N_216), .B(un1_n_s_change_0_1[7]), .Y(
        un1_ten_choice_one_0_1_7));
    NOR2 \dataeight_0_a2[3]  (.A(un1_n_s_change_0_1[3]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_3));
    NOR2A \datafour_0_a2[0]  (.A(N_219), .B(un1_n_s_change_0_1[0]), .Y(
        un1_ten_choice_one_0_3_0));
    NOR2A \dataone_0_a2[10]  (.A(N_222), .B(un1_n_s_change_0_1[10]), 
        .Y(un1_ten_choice_one_0[10]));
    NOR2A \dataseven_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_221), 
        .Y(un1_ten_choice_one_0_6[5]));
    NOR2A \dataone_0_a2[8]  (.A(N_222), .B(un1_n_s_change_0_1[8]), .Y(
        un1_ten_choice_one_0[8]));
    NOR2A \datafour_0_a2[8]  (.A(N_219), .B(un1_n_s_change_0_1[8]), .Y(
        un1_ten_choice_one_0_3_8));
    OR2B \datafive_0_a2_2[0]  (.A(addrout[2]), .B(addrout[0]), .Y(
        N_212));
    NOR2A \datafive_0_a2[0]  (.A(N_217), .B(un1_n_s_change_0_1[0]), .Y(
        un1_ten_choice_one_0_4_0));
    VCC VCC_i (.Y(VCC));
    NOR2A \datafour_0_a2[4]  (.A(N_219), .B(un1_n_s_change_0_1[4]), .Y(
        un1_ten_choice_one_0_3_4));
    NOR2A \dataeight_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_220), 
        .Y(un1_ten_choice_one_0_7_5));
    NOR2 \dataeight_0_a2[11]  (.A(un1_n_s_change_0_1[11]), .B(N_220), 
        .Y(un1_ten_choice_one_0_7_11));
    NOR2 \dataseven_0_a2[4]  (.A(un1_n_s_change_0_1[4]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[4]));
    NOR2A \datafive_0_a2[11]  (.A(N_217), .B(un1_n_s_change_0_1[11]), 
        .Y(un1_ten_choice_one_0_4_11));
    OR2 \datasix_0_a2[7]  (.A(un1_n_s_change_0_1[7]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[7]));
    NOR2 \dataeight_0_a2[7]  (.A(un1_n_s_change_0_1[7]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_7));
    NOR2A \dataone_0_a2[7]  (.A(N_222), .B(un1_n_s_change_0_1[7]), .Y(
        un1_ten_choice_one_0[7]));
    NOR2A \datafour_0_a2[6]  (.A(N_219), .B(un1_n_s_change_0_1[6]), .Y(
        un1_ten_choice_one_0_3_6));
    NOR2A \datatwo_0_a2[6]  (.A(N_216), .B(un1_n_s_change_0_1[6]), .Y(
        un1_ten_choice_one_0_1_6));
    NOR2A \datatwo_0_a2[8]  (.A(N_216), .B(un1_n_s_change_0_1[8]), .Y(
        un1_ten_choice_one_0_1_8));
    NOR2 \datathree_0_a2_0[0]  (.A(N_215), .B(N_210), .Y(N_224));
    NOR2A \datafive_0_a2[7]  (.A(N_217), .B(un1_n_s_change_0_1[7]), .Y(
        un1_ten_choice_one_0_4_7));
    NOR2 \datasix_0_a2[6]  (.A(un1_n_s_change_0_1[6]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[6]));
    NOR2 \dataeight_0_a2[9]  (.A(un1_n_s_change_0_1[9]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_9));
    NOR2 \datasix_0_a2[0]  (.A(un1_n_s_change_0_1[0]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[0]));
    NOR2 \dataseven_0_a2[10]  (.A(un1_n_s_change_0_1[10]), .B(N_221), 
        .Y(un1_ten_choice_one_0_6[10]));
    OR2A \dataone_0_a2[2]  (.A(N_222), .B(un1_n_s_change_0_1[2]), .Y(
        un1_ten_choice_one_0[2]));
    OR2A \datafour_0_a2_1[0]  (.A(addrout[2]), .B(addrout[0]), .Y(
        N_214));
    NOR2 \dataeight_0_a2[10]  (.A(un1_n_s_change_0_1[10]), .B(N_220), 
        .Y(un1_ten_choice_one_0_7_10));
    OR2B \datatwo_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_216), .Y(
        un1_ten_choice_one_0_1_5));
    NOR2 \datafour_0_a2_0[0]  (.A(N_214), .B(N_211), .Y(N_219));
    NOR2A \datafour_0_a2[1]  (.A(N_219), .B(un1_n_s_change_0_1[1]), .Y(
        un1_ten_choice_one_0_3_1));
    NOR2 \datasix_0_a2[10]  (.A(un1_n_s_change_0_1[10]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[10]));
    NOR3 \datathree_0_a2[3]  (.A(N_215), .B(un1_n_s_change_0_1[3]), .C(
        N_210), .Y(un1_ten_choice_one_0_2_2));
    NOR2 \dataeight_0_a2[6]  (.A(un1_n_s_change_0_1[6]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_6));
    NOR2A \datasix_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[5]));
    NOR2B \datafive_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_217), .Y(
        un1_ten_choice_one_0_4_5));
    NOR2 \dataeight_0_a2[8]  (.A(un1_n_s_change_0_1[8]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_8));
    GND GND_i (.Y(GND));
    OR2A \datathree_0_a2[1]  (.A(N_224), .B(un1_n_s_change_0_1[1]), .Y(
        un1_ten_choice_one_0_2_0));
    OR2 \datasix_0_a2[9]  (.A(un1_n_s_change_0_1[9]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[9]));
    OR2A \datafive_0_a2[1]  (.A(N_217), .B(un1_n_s_change_0_1[1]), .Y(
        un1_ten_choice_one_0_4_1));
    NOR2 \datasix_0_a2[8]  (.A(un1_n_s_change_0_1[8]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[8]));
    OR2A \dataone_0_a2_1[0]  (.A(addrout[0]), .B(addrout[2]), .Y(N_215)
        );
    NOR2 \dataone_0_a2_0[0]  (.A(N_215), .B(N_211), .Y(N_222));
    NOR2A \datathree_0_a2[10]  (.A(N_224), .B(un1_n_s_change_0_1[10]), 
        .Y(un1_ten_choice_one_0_2_9));
    OR2 \datasix_0_a2[11]  (.A(un1_n_s_change_0_1[11]), .B(N_223), .Y(
        un1_ten_choice_one_0_5[11]));
    OR2A \dataone_0_a2[9]  (.A(N_222), .B(un1_n_s_change_0_1[9]), .Y(
        un1_ten_choice_one_0[9]));
    OR2 \dataeight_0_a2_0[0]  (.A(dataeight_0_a2_0_0[0]), .B(N_213), 
        .Y(N_220));
    NOR2 \dataseven_0_a2[7]  (.A(un1_n_s_change_0_1[7]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[7]));
    NOR2B \datathree_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_224), 
        .Y(un1_ten_choice_one_0_2_4));
    NOR2 \datafive_0_a2_0[0]  (.A(N_212), .B(N_211), .Y(N_217));
    NOR2A \datafive_0_a2[9]  (.A(N_217), .B(un1_n_s_change_0_1[9]), .Y(
        un1_ten_choice_one_0_4_9));
    OR2A \datatwo_0_a2_1[0]  (.A(addrout[1]), .B(addrout[3]), .Y(N_210)
        );
    NOR2A \datatwo_0_a2[1]  (.A(N_216), .B(un1_n_s_change_0_1[1]), .Y(
        un1_ten_choice_one_0_1_1));
    NOR2 \dataseven_0_a2[6]  (.A(un1_n_s_change_0_1[6]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[6]));
    NOR2A \datatwo_0_a2[2]  (.A(N_216), .B(un1_n_s_change_0_1[2]), .Y(
        un1_ten_choice_one_0_1_2));
    NOR2A \datafive_0_a2[4]  (.A(N_217), .B(un1_n_s_change_0_1[4]), .Y(
        un1_ten_choice_one_0_4_4));
    NOR2A \datatwo_0_a2[0]  (.A(N_216), .B(un1_n_s_change_0_1[0]), .Y(
        un1_ten_choice_one_0_1_0));
    NOR2 \dataeight_0_a2[0]  (.A(un1_n_s_change_0_1[0]), .B(N_220), .Y(
        un1_ten_choice_one_0_7_0));
    OR2A \dataeight_0_a2_0_0[0]  (.A(addrout[3]), .B(addrout[1]), .Y(
        dataeight_0_a2_0_0[0]));
    NOR2A \datafour_0_a2[3]  (.A(N_219), .B(un1_n_s_change_0_1[3]), .Y(
        un1_ten_choice_one_0_3_3));
    NOR2A \datathree_0_a2[4]  (.A(N_224), .B(un1_n_s_change_0_1[4]), 
        .Y(un1_ten_choice_one_0_2_3));
    NOR2A \datafour_0_a2[7]  (.A(N_219), .B(un1_n_s_change_0_1[7]), .Y(
        un1_ten_choice_one_0_3_7));
    NOR2A \datafour_0_a2[11]  (.A(N_219), .B(un1_n_s_change_0_1[11]), 
        .Y(un1_ten_choice_one_0_3_11));
    NOR2A \datathree_0_a2[11]  (.A(N_224), .B(un1_n_s_change_0_1[11]), 
        .Y(un1_ten_choice_one_0_2_10));
    NOR2A \datafour_0_a2[10]  (.A(N_219), .B(un1_n_s_change_0_1[10]), 
        .Y(un1_ten_choice_one_0_3_10));
    NOR2 \dataseven_0_a2[8]  (.A(un1_n_s_change_0_1[8]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[8]));
    NOR2 \datatwo_0_a2_0[0]  (.A(N_213), .B(N_210), .Y(N_216));
    NOR2A \datathree_0_a2[9]  (.A(N_224), .B(un1_n_s_change_0_1[9]), 
        .Y(un1_ten_choice_one_0_2_8));
    NOR2A \datathree_0_a2[7]  (.A(N_224), .B(un1_n_s_change_0_1[7]), 
        .Y(un1_ten_choice_one_0_2_6));
    NOR2A \dataone_0_a2[11]  (.A(N_222), .B(un1_n_s_change_0_1[11]), 
        .Y(un1_ten_choice_one_0[11]));
    NOR2 \dataseven_0_a2[9]  (.A(un1_n_s_change_0_1[9]), .B(N_221), .Y(
        un1_ten_choice_one_0_6[9]));
    NOR2A \datafour_0_a2[9]  (.A(N_219), .B(un1_n_s_change_0_1[9]), .Y(
        un1_ten_choice_one_0_3_9));
    OR2 \datafive_0_a2_1[0]  (.A(addrout[3]), .B(addrout[1]), .Y(N_211)
        );
    NOR2B \datafour_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_219), .Y(
        un1_ten_choice_one_0_3_5));
    NOR2A \datatwo_0_a2[4]  (.A(N_216), .B(un1_n_s_change_0_1[4]), .Y(
        un1_ten_choice_one_0_1_4));
    NOR2A \datathree_0_a2[6]  (.A(N_224), .B(un1_n_s_change_0_1[6]), 
        .Y(un1_ten_choice_one_0_2_5));
    NOR2A \dataone_0_a2[4]  (.A(N_222), .B(un1_n_s_change_0_1[4]), .Y(
        un1_ten_choice_one_0[4]));
    NOR2A \dataone_0_a2[6]  (.A(N_222), .B(un1_n_s_change_0_1[6]), .Y(
        un1_ten_choice_one_0[6]));
    NOR2A \dataone_0_a2[1]  (.A(N_222), .B(un1_n_s_change_0_1[1]), .Y(
        un1_ten_choice_one_0[1]));
    NOR2A \datafive_0_a2[6]  (.A(N_217), .B(un1_n_s_change_0_1[6]), .Y(
        un1_ten_choice_one_0_4_6));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR2A \datatwo_0_a2[11]  (.A(N_216), .B(un1_n_s_change_0_1[11]), 
        .Y(un1_ten_choice_one_0_1_11));
    NOR2B \dataone_0_a2[5]  (.A(un1_n_s_change_0_1[5]), .B(N_222), .Y(
        un1_ten_choice_one_0[5]));
    
endmodule


module add_reg_add_reg_2_7(
       addresult_RNIVJME,
       signal_data_0_iv_i_2,
       signal_data_iv_0_0_3,
       signal_data_iv_0_3_0,
       signal_data_iv_0_3_3,
       signal_data_iv_0_3_2,
       ADC_c,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_4_0,
       un1_ten_choice_one_0_4_3,
       un1_ten_choice_one_0_4_1,
       un1_ten_choice_one_0_4_4,
       un1_ten_choice_one_0_4_5,
       un1_ten_choice_one_0_4_7,
       un1_ten_choice_one_0_4_8,
       un1_ten_choice_one_0_4_9,
       un1_ten_choice_one_0_4_10,
       un1_ten_choice_one_0_4_11,
       un1_ten_choice_one_0_4_6,
       un1_add_reg_4_i_2,
       un1_add_reg_4_i_0,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_218,
       N_186,
       N_88,
       N_104,
       N_249,
       N_202,
       N_250,
       N_249_0,
       N_235,
       N_212,
       N_211,
       N_188,
       N_177,
       N_145,
       N_137,
       N_129,
       N_121,
       N_153,
       N_169,
       N_253,
       N_237,
       N_204,
       N_220,
       N_263,
       top_code_0_n_s_ctrl_0,
       N_217
    );
input  [4:4] addresult_RNIVJME;
output [11:4] signal_data_0_iv_i_2;
output [1:1] signal_data_iv_0_0_3;
output signal_data_iv_0_3_0;
output signal_data_iv_0_3_3;
output signal_data_iv_0_3_2;
input  [2:0] ADC_c;
input  [3:2] un1_n_s_change_0_1;
input  un1_ten_choice_one_0_4_0;
input  un1_ten_choice_one_0_4_3;
input  un1_ten_choice_one_0_4_1;
input  un1_ten_choice_one_0_4_4;
input  un1_ten_choice_one_0_4_5;
input  un1_ten_choice_one_0_4_7;
input  un1_ten_choice_one_0_4_8;
input  un1_ten_choice_one_0_4_9;
input  un1_ten_choice_one_0_4_10;
input  un1_ten_choice_one_0_4_11;
input  un1_ten_choice_one_0_4_6;
output un1_add_reg_4_i_2;
output un1_add_reg_4_i_0;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
output N_218;
output N_186;
output N_88;
output N_104;
input  N_249;
output N_202;
input  N_250;
input  N_249_0;
output N_235;
input  N_212;
input  N_211;
input  N_188;
input  N_177;
input  N_145;
input  N_137;
input  N_129;
input  N_121;
input  N_153;
input  N_169;
input  N_253;
input  N_237;
input  N_204;
input  N_220;
input  N_263;
input  top_code_0_n_s_ctrl_0;
input  N_217;

    wire ADD_20x20_slow_I13_CO1_0, \addresult_2[12] , 
        ADD_20x20_slow_I6_S_0_0, \addresult_2[6] , 
        ADD_20x20_slow_I2_S_0_0, \addresult_2[2] , 
        ADD_20x20_slow_I5_CO1_0_tz_0, \addresult_2[4] , N232, 
        \addresult_2[5] , ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_1, 
        ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0, 
        ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0, 
        ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_0, 
        ADD_20x20_slow_I2_un1_CO1_N_15, \addresult_2[3] , 
        \addresult_2[1] , \addresult_2[11] , \addresult_1[7] , 
        \addresult_2[8] , \addresult_2[9] , \addresult_2[10] , 
        \addresult_2[0] , \un3_addresult[11] , I10_un1_CO1, 
        \un3_addresult[10] , N244, \un3_addresult[9] , I8_un1_CO1, 
        \un3_addresult[8] , N240, \un3_addresult[7] , I6_un1_CO1, 
        \un3_addresult[6] , N236, \un3_addresult[5] , I4_un1_CO1, 
        \un3_addresult[4] , \un3_addresult[2] , 
        ADD_20x20_slow_I1_CO1_0, I1_un3_CO1, \un3_addresult[1] , 
        I0_un1_CO1, \un3_addresult[3] , I2_un1_CO1_i, 
        ADD_20x20_slow_I3_CO1_0, I3_un2_CO1_i, 
        ADD_20x20_slow_I2_un1_CO1tt_m1_e, ADD_20x20_slow_I5_CO1_0, 
        ADD_20x20_slow_I4_un1_CO1_0, I5_un5_CO1, N248, I14_un1_CO1, 
        \addresult_2[14] , I16_un1_CO1, \addresult_2[16] , 
        \un3_addresult[14] , \un3_addresult[15] , \un3_addresult[16] , 
        \un3_addresult[17] , \addresult_2[17] , \un3_addresult[13] , 
        \un3_addresult[12] , \addresult_2[19] , \un3_addresult[0] , 
        \addresult_2[18] , \un3_addresult[19] , N270, 
        \un3_addresult[18] , GND, VCC, GND_0, VCC_0;
    
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        un1_ten_choice_one_0_4_11), .B(\addresult_2[11] ), .C(
        I10_un1_CO1), .Y(\un3_addresult[11] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[12] ));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_4_8), .B(\addresult_2[8] ), .C(N240), .Y(
        \un3_addresult[8] ));
    AOI1B \addresult_RNIG75R[0]  (.A(\addresult_2[0] ), .B(N_263), .C(
        N_188), .Y(signal_data_iv_0_3_0));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[10] ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[6] ));
    OR2B un3_addresult_ADD_20x20_slow_I3_CO1 (.A(I3_un2_CO1_i), .B(
        ADD_20x20_slow_I3_CO1_0), .Y(N232));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[8] ));
    OA1 \addresult_RNIPQMP[5]  (.A(N_253), .B(\addresult_2[5] ), .C(
        N_169), .Y(signal_data_0_iv_i_2[5]));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(
        un1_ten_choice_one_0_4_1), .B(\addresult_2[1] ), .C(I0_un1_CO1)
        , .Y(\un3_addresult[1] ));
    OR2A un3_addresult_ADD_20x20_slow_I1_un3_CO1 (.A(ADC_c[1]), .B(
        I0_un1_CO1), .Y(I1_un3_CO1));
    OR3A \addresult_RNIJ70G[16]  (.A(\addresult_2[16] ), .B(N_249), .C(
        N_250), .Y(N_186));
    DFN1P0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        un1_add_reg_4_i_2));
    VCC VCC_i (.Y(VCC));
    OAI1 un3_addresult_ADD_20x20_slow_I5_CO1_0 (.A(
        ADD_20x20_slow_I4_un1_CO1_0), .B(ADD_20x20_slow_I5_CO1_0_tz_0), 
        .C(un1_ten_choice_one_0_4_5), .Y(ADD_20x20_slow_I5_CO1_0));
    NOR2B un3_addresult_ADD_20x20_slow_I2_un1_CO1tt_m1_e (.A(
        \addresult_2[0] ), .B(ADC_c[0]), .Y(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e));
    MAJ3 un3_addresult_ADD_20x20_slow_I11_CO1 (.A(I10_un1_CO1), .B(
        \addresult_2[11] ), .C(un1_ten_choice_one_0_4_11), .Y(N248));
    OR2B un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I5_un5_CO1), .B(
        ADD_20x20_slow_I5_CO1_0), .Y(N236));
    AOI1B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_1 (.A(
        ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0), .B(
        ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0), .C(
        ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_0), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_1));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[4] ));
    OR2A un3_addresult_ADD_20x20_slow_I3_un2_CO1 (.A(\addresult_2[3] ), 
        .B(un1_ten_choice_one_0_4_3), .Y(I3_un2_CO1_i));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0_4_0), .B(\addresult_2[0] ), .Y(
        \un3_addresult[0] ));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[16] ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_4_5), .B(\addresult_2[5] ), .C(I4_un1_CO1)
        , .Y(\un3_addresult[5] ));
    OR2 \addresult_RNITTFB[14]  (.A(\addresult_2[14] ), .B(N_253), .Y(
        N_104));
    OAI1 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0 (.A(
        ADC_c[1]), .B(ADD_20x20_slow_I2_un1_CO1tt_m1_e), .C(
        \addresult_2[1] ), .Y(ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0));
    AX1 un3_addresult_ADD_20x20_slow_I14_S_0 (.A(
        ADD_20x20_slow_I13_CO1_0), .B(N248), .C(\addresult_2[14] ), .Y(
        \un3_addresult[14] ));
    XOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0_4_4), .B(\addresult_2[4] ), .C(N232), .Y(
        \un3_addresult[4] ));
    XOR2 un3_addresult_ADD_20x20_slow_I18_S_0 (.A(\addresult_2[18] ), 
        .B(N270), .Y(\un3_addresult[18] ));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[5] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_2[8] ), .C(un1_ten_choice_one_0_4_8), .Y(I8_un1_CO1)
        );
    OR2B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_a3_1 (.A(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e), .B(ADC_c[1]), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_15));
    AX1C un3_addresult_ADD_20x20_slow_I19_Y_0 (.A(N270), .B(
        \addresult_2[18] ), .C(\addresult_2[19] ), .Y(
        \un3_addresult[19] ));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[2] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult_1[7] ), .C(un1_ten_choice_one_0_4_7), .Y(N240));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0_0 (.A(\addresult_2[6] ), 
        .B(un1_ten_choice_one_0_4_6), .Y(ADD_20x20_slow_I6_S_0_0));
    OR3B un3_addresult_ADD_20x20_slow_I14_un1_CO1 (.A(N248), .B(
        \addresult_2[14] ), .C(ADD_20x20_slow_I13_CO1_0), .Y(
        I14_un1_CO1));
    OA1 \addresult_RNI1RNP[9]  (.A(N_253), .B(\addresult_2[9] ), .C(
        N_137), .Y(signal_data_0_iv_i_2[9]));
    OR2B un3_addresult_ADD_20x20_slow_I5_un5_CO1 (.A(\addresult_2[5] ), 
        .B(I4_un1_CO1), .Y(I5_un5_CO1));
    AX1B un3_addresult_ADD_20x20_slow_I16_S_0 (.A(I14_un1_CO1), .B(
        un1_add_reg_4_i_2), .C(\addresult_2[16] ), .Y(
        \un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[3] ));
    OA1 \addresult_RNITANP[7]  (.A(N_253), .B(\addresult_1[7] ), .C(
        N_121), .Y(signal_data_0_iv_i_2[7]));
    XNOR2 un3_addresult_ADD_20x20_slow_I17_S_0 (.A(\addresult_2[17] ), 
        .B(I16_un1_CO1), .Y(\un3_addresult[17] ));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[14] ));
    AO1B un3_addresult_ADD_20x20_slow_I1_CO1_0 (.A(
        un1_ten_choice_one_0_4_1), .B(I0_un1_CO1), .C(\addresult_2[1] )
        , .Y(ADD_20x20_slow_I1_CO1_0));
    XOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(\addresult_2[12] ), 
        .B(N248), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    AO1 un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(\addresult_2[4] ), 
        .B(N232), .C(ADD_20x20_slow_I4_un1_CO1_0), .Y(I4_un1_CO1));
    OA1B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_0 (.A(
        ADC_c[2]), .B(\addresult_2[2] ), .C(top_code_0_n_s_ctrl_0), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_0));
    OR3A un3_addresult_ADD_20x20_slow_I16_un1_CO1 (.A(
        \addresult_2[16] ), .B(I14_un1_CO1), .C(un1_add_reg_4_i_2), .Y(
        I16_un1_CO1));
    OR2 \addresult_RNIRTFB[12]  (.A(\addresult_2[12] ), .B(N_253), .Y(
        N_88));
    AOI1B \addresult_RNIIB5R[1]  (.A(\addresult_2[1] ), .B(N_263), .C(
        N_237), .Y(signal_data_iv_0_0_3[1]));
    NOR2A un3_addresult_ADD_20x20_slow_I17_CO1 (.A(\addresult_2[17] ), 
        .B(I16_un1_CO1), .Y(N270));
    OR3A \addresult_RNIK70G[17]  (.A(\addresult_2[17] ), .B(N_249_0), 
        .C(N_250), .Y(N_235));
    XNOR2 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(un1_add_reg_4_i_2), 
        .B(I14_un1_CO1), .Y(\un3_addresult[15] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult_2[10] ), .C(un1_ten_choice_one_0_4_10), .Y(
        I10_un1_CO1));
    OA1 \addresult_RNI93LI[11]  (.A(N_253), .B(\addresult_2[11] ), .C(
        N_153), .Y(signal_data_0_iv_i_2[11]));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[11] ));
    OA1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0 (.A(N232), .B(
        \addresult_2[4] ), .C(un1_ten_choice_one_0_4_4), .Y(
        ADD_20x20_slow_I4_un1_CO1_0));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[17] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1), .B(
        \addresult_2[9] ), .C(un1_ten_choice_one_0_4_9), .Y(N244));
    AO1 un3_addresult_ADD_20x20_slow_I5_CO1_0_tz_0 (.A(
        \addresult_2[4] ), .B(N232), .C(\addresult_2[5] ), .Y(
        ADD_20x20_slow_I5_CO1_0_tz_0));
    AX1A un3_addresult_ADD_20x20_slow_I2_S_0_0 (.A(
        un1_n_s_change_0_1[2]), .B(N_217), .C(\addresult_2[2] ), .Y(
        ADD_20x20_slow_I2_S_0_0));
    OR2A un3_addresult_ADD_20x20_slow_I13_CO1_0 (.A(\addresult_2[12] ), 
        .B(un1_add_reg_4_i_0), .Y(ADD_20x20_slow_I13_CO1_0));
    MAJ3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult_2[6] ), .C(un1_ten_choice_one_0_4_6), .Y(I6_un1_CO1)
        );
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_4_10), .B(\addresult_2[10] ), .C(N244), 
        .Y(\un3_addresult[10] ));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_1[7] ));
    AX1C un3_addresult_ADD_20x20_slow_I13_S_0 (.A(N248), .B(
        \addresult_2[12] ), .C(un1_add_reg_4_i_0), .Y(
        \un3_addresult[13] ));
    XOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(I2_un1_CO1_i), .B(
        \addresult_2[3] ), .C(un1_ten_choice_one_0_4_3), .Y(
        \un3_addresult[3] ));
    OA1 \addresult_RNIR2NP[6]  (.A(N_253), .B(\addresult_2[6] ), .C(
        N_177), .Y(signal_data_0_iv_i_2[6]));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[18] ));
    OR3A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e (.A(
        ADD_20x20_slow_I2_un1_CO1_m11_i_m2_e_1), .B(N_211), .C(N_212), 
        .Y(I2_un1_CO1_i));
    AOI1B \addresult_RNIMJ5R[3]  (.A(\addresult_2[3] ), .B(N_263), .C(
        N_204), .Y(signal_data_iv_0_3_3));
    OA1 \addresult_RNINIMP[4]  (.A(N_253), .B(\addresult_2[4] ), .C(
        addresult_RNIVJME[4]), .Y(signal_data_0_iv_i_2[4]));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        ADD_20x20_slow_I6_S_0_0), .B(N236), .Y(\un3_addresult[6] ));
    AOI1B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0_0 (.A(
        \addresult_2[2] ), .B(ADC_c[2]), .C(
        ADD_20x20_slow_I2_un1_CO1_N_15), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0));
    OA1 \addresult_RNI73LI[10]  (.A(N_253), .B(\addresult_2[10] ), .C(
        N_145), .Y(signal_data_0_iv_i_2[10]));
    DFN1P0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        un1_add_reg_4_i_0));
    OR3A \addresult_RNIM70G[19]  (.A(\addresult_2[19] ), .B(N_249), .C(
        N_250), .Y(N_202));
    AOI1B \addresult_RNIKF5R[2]  (.A(\addresult_2[2] ), .B(N_263), .C(
        N_220), .Y(signal_data_iv_0_3_2));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[9] ));
    DFN1C0 \addresult[19]  (.D(\un3_addresult[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[19] ));
    AO1A un3_addresult_ADD_20x20_slow_I3_CO1_0 (.A(\addresult_2[3] ), 
        .B(un1_n_s_change_0_1[3]), .C(I2_un1_CO1_i), .Y(
        ADD_20x20_slow_I3_CO1_0));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[0] ));
    OR2B un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(
        un1_ten_choice_one_0_4_0), .B(\addresult_2[0] ), .Y(I0_un1_CO1)
        );
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0_4_7), .B(\addresult_1[7] ), .C(I6_un1_CO1)
        , .Y(\un3_addresult[7] ));
    OR3A \addresult_RNIL70G[18]  (.A(\addresult_2[18] ), .B(N_249), .C(
        N_250), .Y(N_218));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_4_9), .B(\addresult_2[9] ), .C(I8_un1_CO1)
        , .Y(\un3_addresult[9] ));
    AX1C un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        ADD_20x20_slow_I1_CO1_0), .B(I1_un3_CO1), .C(
        ADD_20x20_slow_I2_S_0_0), .Y(\un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    OA1 \addresult_RNIVINP[8]  (.A(N_253), .B(\addresult_2[8] ), .C(
        N_129), .Y(signal_data_0_iv_i_2[8]));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[1] ));
    
endmodule


module s_clk_div4(
       s_acq_change_0_s_rst,
       ddsclkout_c,
       clkout,
       scan_scale_sw_0_s_start,
       signalclkctrl_0_entop
    );
input  s_acq_change_0_s_rst;
input  ddsclkout_c;
output clkout;
input  scan_scale_sw_0_s_start;
input  signalclkctrl_0_entop;

    wire clkout_1_sqmuxa, count_net_1, clkout_4, count_RNO_net_1, GND, 
        VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 count (.D(count_RNO_net_1), .CLK(ddsclkout_c), .CLR(
        s_acq_change_0_s_rst), .Q(count_net_1));
    NOR3B clkout_RNO (.A(signalclkctrl_0_entop), .B(
        scan_scale_sw_0_s_start), .C(clkout), .Y(clkout_4));
    DFN1E0C0 clkout_inst_1 (.D(clkout_4), .CLK(ddsclkout_c), .CLR(
        s_acq_change_0_s_rst), .E(clkout_1_sqmuxa), .Q(clkout));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    AX1C count_RNO (.A(signalclkctrl_0_entop), .B(
        scan_scale_sw_0_s_start), .C(count_net_1), .Y(count_RNO_net_1));
    NOR3B clkout_RNO_0 (.A(signalclkctrl_0_entop), .B(
        scan_scale_sw_0_s_start), .C(count_net_1), .Y(clkout_1_sqmuxa));
    
endmodule


module ctrl_addr(
       s_periodnum,
       addrout,
       s_acq_change_0_s_load_0,
       GLA,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add
    );
input  [3:0] s_periodnum;
output [3:0] addrout;
input  s_acq_change_0_s_load_0;
input  GLA;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;

    wire N_7, \addrout_RNI1LRG[1]_net_1 , \addrout_RNI0HRG[0]_net_1 , 
        addrout14_NE_1, \datareg[3]_net_1 , addrout14_0_i, 
        addrout14_NE_0, \datareg[1]_net_1 , addrout14_2_i, 
        \addrout_RNI2PRG[2]_net_1 , \addrout_RNI3TRG[3]_net_1 , 
        \datareg[0]_net_1 , \datareg[2]_net_1 , \addrout_3[0] , 
        \addrout_3[1] , \addrout_3[2] , \addrout_3[3] , N_4, GND, VCC, 
        GND_0, VCC_0;
    
    DFN1E1 \datareg[2]  (.D(s_periodnum[2]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\datareg[2]_net_1 ));
    AOI1B \addrout_RNI1LRG[1]  (.A(addrout14_NE_1), .B(addrout14_NE_0), 
        .C(addrout[1]), .Y(\addrout_RNI1LRG[1]_net_1 ));
    AOI1B \addrout_RNI2PRG[2]  (.A(addrout14_NE_1), .B(addrout14_NE_0), 
        .C(addrout[2]), .Y(\addrout_RNI2PRG[2]_net_1 ));
    NOR2B addrout_3_I_8 (.A(\addrout_RNI1LRG[1]_net_1 ), .B(
        \addrout_RNI0HRG[0]_net_1 ), .Y(N_7));
    XOR2 addrout_3_I_13 (.A(N_4), .B(\addrout_RNI3TRG[3]_net_1 ), .Y(
        \addrout_3[3] ));
    GND GND_i_0 (.Y(GND_0));
    DFN0C0 \addrout[2]  (.D(\addrout_3[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addrout[2]));
    VCC VCC_i (.Y(VCC));
    AOI1B \addrout_RNI0HRG[0]  (.A(addrout14_NE_1), .B(addrout14_NE_0), 
        .C(addrout[0]), .Y(\addrout_RNI0HRG[0]_net_1 ));
    DFN1E1 \datareg[1]  (.D(s_periodnum[1]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\datareg[1]_net_1 ));
    AND3 addrout_3_I_12 (.A(\addrout_RNI0HRG[0]_net_1 ), .B(
        \addrout_RNI1LRG[1]_net_1 ), .C(\addrout_RNI2PRG[2]_net_1 ), 
        .Y(N_4));
    XNOR2 \datareg_RNI7S54[2]  (.A(addrout[2]), .B(\datareg[2]_net_1 ), 
        .Y(addrout14_2_i));
    GND GND_i (.Y(GND));
    AOI1B \addrout_RNI3TRG[3]  (.A(addrout14_NE_1), .B(addrout14_NE_0), 
        .C(addrout[3]), .Y(\addrout_RNI3TRG[3]_net_1 ));
    DFN1E1 \datareg[0]  (.D(s_periodnum[0]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\datareg[0]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    XA1A \datareg_RNICGB8[3]  (.A(\datareg[3]_net_1 ), .B(addrout[3]), 
        .C(addrout14_0_i), .Y(addrout14_NE_1));
    XOR2 addrout_3_I_5 (.A(\addrout_RNI0HRG[0]_net_1 ), .B(
        \addrout_RNI1LRG[1]_net_1 ), .Y(\addrout_3[1] ));
    DFN0C0 \addrout[1]  (.D(\addrout_3[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addrout[1]));
    DFN0P0 \addrout[0]  (.D(\addrout_3[0] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        addrout[0]));
    DFN0C0 \addrout[3]  (.D(\addrout_3[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addrout[3]));
    DFN1E1 \datareg[3]  (.D(s_periodnum[3]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\datareg[3]_net_1 ));
    XOR2 addrout_3_I_9 (.A(N_7), .B(\addrout_RNI2PRG[2]_net_1 ), .Y(
        \addrout_3[2] ));
    XA1A \datareg_RNICGB8[1]  (.A(\datareg[1]_net_1 ), .B(addrout[1]), 
        .C(addrout14_2_i), .Y(addrout14_NE_0));
    INV addrout_3_I_4 (.A(\addrout_RNI0HRG[0]_net_1 ), .Y(
        \addrout_3[0] ));
    XNOR2 \datareg_RNI3C54[0]  (.A(addrout[0]), .B(\datareg[0]_net_1 ), 
        .Y(addrout14_0_i));
    
endmodule


module add_reg_add_reg_2_3(
       addresult_RNIDU3E,
       signal_data_iv_0_0_6,
       signal_data_iv_0_6_0,
       signal_data_iv_0_6_3,
       signal_data_iv_0_6_2,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_1_0,
       un1_ten_choice_one_0_1_2,
       un1_ten_choice_one_0_1_10,
       un1_ten_choice_one_0_1_5,
       un1_ten_choice_one_0_1_9,
       un1_ten_choice_one_0_1_7,
       un1_ten_choice_one_0_1_1,
       un1_ten_choice_one_0_1_8,
       un1_ten_choice_one_0_1_4,
       un1_ten_choice_one_0_1_6,
       un1_ten_choice_one_0_1_11,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_249,
       N_224,
       N_91,
       N_107,
       N_192,
       N_208,
       N_251,
       N_249_0,
       N_241,
       N_179,
       N_171,
       N_155,
       N_147,
       N_139,
       N_131,
       N_123,
       N_115,
       N_254,
       N_99,
       N_194,
       N_243,
       N_210_0,
       N_226,
       N_273,
       N_213,
       N_210,
       N_216
    );
output [4:4] addresult_RNIDU3E;
output [1:1] signal_data_iv_0_0_6;
output signal_data_iv_0_6_0;
output signal_data_iv_0_6_3;
output signal_data_iv_0_6_2;
input  [3:0] un1_n_s_change_0_1;
input  un1_ten_choice_one_0_1_0;
input  un1_ten_choice_one_0_1_2;
input  un1_ten_choice_one_0_1_10;
input  un1_ten_choice_one_0_1_5;
input  un1_ten_choice_one_0_1_9;
input  un1_ten_choice_one_0_1_7;
input  un1_ten_choice_one_0_1_1;
input  un1_ten_choice_one_0_1_8;
input  un1_ten_choice_one_0_1_4;
input  un1_ten_choice_one_0_1_6;
input  un1_ten_choice_one_0_1_11;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
input  N_249;
output N_224;
output N_91;
output N_107;
output N_192;
output N_208;
input  N_251;
input  N_249_0;
output N_241;
output N_179;
output N_171;
output N_155;
output N_147;
output N_139;
output N_131;
output N_123;
output N_115;
input  N_254;
output N_99;
input  N_194;
input  N_243;
input  N_210_0;
input  N_226;
input  N_273;
input  N_213;
input  N_210;
input  N_216;

    wire ADD_20x20_slow_I11_S_0_0, \addresult_4[11] , 
        ADD_20x20_slow_I10_un1_CO1_0_tz_0, \addresult_4[9] , 
        I8_un1_CO1, \addresult_4[10] , ADD_20x20_slow_I6_S_0_0, 
        \addresult_4[6] , ADD_20x20_slow_I3_S_0_0, \addresult_4[3] , 
        ADD_20x20_slow_I4_S_0_0, \addresult_4[4] , 
        ADD_20x20_slow_I8_un1_CO1_0_m6_0, \addresult_4[8] , 
        ADD_20x20_slow_I1_S_0_0, \addresult_4[1] , 
        ADD_20x20_slow_I3_CO1_m12_0_1, 
        ADD_20x20_slow_I3_CO1_m12_0_a5_0_1, 
        ADD_20x20_slow_I3_CO1tt_m1_0_a2, 
        ADD_20x20_slow_I3_CO1_m12_0_a5, ADD_20x20_slow_I3_CO1_m12_0_0, 
        ADD_20x20_slow_I3_CO1_N_16, ADD_20x20_slow_I1_CO1_0, 
        ADD_20x20_slow_I1_un3_CO1_m2_0_a2_2, 
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_2, 
        ADD_20x20_slow_I3_CO1_m3_e, ADD_20x20_slow_I3_CO1_m12_0_o5, 
        ADD_20x20_slow_I3_CO1_m12_0_o5_0, \addresult_4[0] , 
        ADD_20x20_slow_I1_un3_CO1_m2_0_a2_0, 
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_0, 
        ADD_20x20_slow_I19_Y_0_m6_e_3, \addresult_4[12] , 
        \addresult_4[18] , \addresult_4[17] , 
        ADD_20x20_slow_I19_Y_0_m6_e_2, \addresult_3[15] , 
        \addresult_4[16] , ADD_20x20_slow_I19_Y_0_m6_e_1, 
        \addresult_3[13] , \addresult_4[14] , \addresult_4[2] , 
        \addresult_RNIM85T1[7]_net_1 , d_N_8_2, d_N_7_2, 
        \addresult_3[7] , \addresult_RNI1O4G[7]_net_1 , 
        ADD_20x20_slow_I8_un1_CO1_0_N_7_i, ADD_20x20_slow_I7_S_0_0, 
        \un3_addresult[11] , I10_un1_CO1, \un3_addresult[9] , 
        \un3_addresult[6] , N236, \un3_addresult[5] , 
        \un1_add_reg_1_i[5] , I4_un1_CO1_i, \un3_addresult[4] , 
        ADD_20x20_slow_I3_CO1_m12_0, \un3_addresult[3] , 
        ADD_20x20_slow_I2_un1_CO1_0, I2_un4_CO1, \un3_addresult[10] , 
        N244, \un3_addresult[8] , N240, N228, \un3_addresult[2] , 
        \un3_addresult[1] , ADD_20x20_slow_I19_Y_0_m6_e_2_0, 
        ADD_20x20_slow_I3_CO1_N_9, \un3_addresult[7] , I6_un1_CO1, 
        ADD_20x20_slow_I8_un1_CO1_0, r_N_2_1_i_0, 
        \addresult_RNO_2[19] , r_N_7_i, \addresult_4[19] , 
        ADD_20x20_slow_I10_un1_CO1_0, ADD_20x20_slow_I9_CO1_0, 
        I10_un5_CO1, N254, N262, \un3_addresult[12] , 
        \un3_addresult[13] , \un3_addresult[14] , \un3_addresult[15] , 
        \un3_addresult[16] , \un3_addresult[18] , N270, 
        \un3_addresult[17] , \un3_addresult[0] , GND, VCC, GND_0, 
        VCC_0;
    
    XOR2 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        ADD_20x20_slow_I11_S_0_0), .B(I10_un1_CO1), .Y(
        \un3_addresult[11] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[12] ));
    OR2 \addresult_RNIDU3E[4]  (.A(\addresult_4[4] ), .B(N_254), .Y(
        addresult_RNIDU3E[4]));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_1_8), .B(\addresult_4[8] ), .C(N240), .Y(
        \un3_addresult[8] ));
    OR2 \addresult_RNIRKFE[13]  (.A(\addresult_3[13] ), .B(N_254), .Y(
        N_99));
    MIN3 \addresult_RNIEPOJ42[11]  (.A(I10_un1_CO1), .B(
        \addresult_4[11] ), .C(un1_ten_choice_one_0_1_11), .Y(r_N_7_i));
    OR2A un3_addresult_ADD_20x20_slow_I2_un4_CO1 (.A(N228), .B(
        un1_n_s_change_0_1[2]), .Y(I2_un4_CO1));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[10] ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[6] ));
    OR2 \addresult_RNISKFE[14]  (.A(\addresult_4[14] ), .B(N_254), .Y(
        N_107));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[8] ));
    AX1A un3_addresult_ADD_20x20_slow_I3_S_0_0 (.A(
        un1_n_s_change_0_1[3]), .B(N_216), .C(\addresult_4[3] ), .Y(
        ADD_20x20_slow_I3_S_0_0));
    XOR2 un3_addresult_ADD_20x20_slow_I4_S_0_0 (.A(\addresult_4[4] ), 
        .B(un1_ten_choice_one_0_1_4), .Y(ADD_20x20_slow_I4_S_0_0));
    OR3 \addresult_RNI2G901[8]  (.A(un1_ten_choice_one_0_1_6), .B(
        \addresult_4[8] ), .C(\addresult_RNI1O4G[7]_net_1 ), .Y(
        d_N_7_2));
    NOR3B un3_addresult_ADD_20x20_slow_I1_un3_CO1_m2_0_a2_2 (.A(
        \addresult_4[0] ), .B(ADD_20x20_slow_I1_un3_CO1_m2_0_a2_0), .C(
        N_213), .Y(ADD_20x20_slow_I1_un3_CO1_m2_0_a2_2));
    AX1C un3_addresult_ADD_20x20_slow_I1_S_0 (.A(\addresult_4[0] ), .B(
        un1_ten_choice_one_0_1_0), .C(ADD_20x20_slow_I1_S_0_0), .Y(
        \un3_addresult[1] ));
    NOR2 un3_addresult_ADD_20x20_slow_I3_CO1_m12_0 (.A(
        ADD_20x20_slow_I3_CO1_m12_0_1), .B(
        ADD_20x20_slow_I3_CO1_m12_0_0), .Y(ADD_20x20_slow_I3_CO1_m12_0)
        );
    OR2 \addresult_RNIGA4E[7]  (.A(\addresult_3[7] ), .B(N_254), .Y(
        N_123));
    NOR2B un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_o5_1 (.A(N_216), 
        .B(ADD_20x20_slow_I3_CO1_m12_0_o5), .Y(
        ADD_20x20_slow_I3_CO1_N_9));
    AOI1B \addresult_RNI4U811[0]  (.A(\addresult_4[0] ), .B(N_273), .C(
        N_194), .Y(signal_data_iv_0_6_0));
    NOR2 un3_addresult_ADD_20x20_slow_I1_un3_CO1_m2_0_a2_0 (.A(
        un1_n_s_change_0_1[0]), .B(un1_n_s_change_0_1[1]), .Y(
        ADD_20x20_slow_I1_un3_CO1_m2_0_a2_0));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[15] ));
    XNOR2 \addresult_RNO[19]  (.A(r_N_7_i), .B(\addresult_4[19] ), .Y(
        \addresult_RNO_2[19] ));
    NOR2B \addresult_RNI1O4G[7]  (.A(un1_ten_choice_one_0_1_7), .B(
        \addresult_3[7] ), .Y(\addresult_RNI1O4G[7]_net_1 ));
    VCC VCC_i (.Y(VCC));
    MIN3 un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I4_un1_CO1_i), .B(
        \un1_add_reg_1_i[5] ), .C(un1_ten_choice_one_0_1_5), .Y(N236));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[4] ));
    AO1D un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_1 (.A(
        ADD_20x20_slow_I3_CO1_m12_0_a5_0_1), .B(
        ADD_20x20_slow_I3_CO1tt_m1_0_a2), .C(
        ADD_20x20_slow_I3_CO1_m12_0_a5), .Y(
        ADD_20x20_slow_I3_CO1_m12_0_1));
    OR3B un3_addresult_ADD_20x20_slow_I15_CO1 (.A(\addresult_4[14] ), 
        .B(\addresult_3[15] ), .C(N254), .Y(N262));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0_1_0), .B(\addresult_4[0] ), .Y(
        \un3_addresult[0] ));
    OR2 \addresult_RNIOKFE[10]  (.A(\addresult_4[10] ), .B(N_254), .Y(
        N_147));
    OR3B un3_addresult_ADD_20x20_slow_I13_CO1 (.A(\addresult_4[12] ), 
        .B(\addresult_3[13] ), .C(r_N_7_i), .Y(N254));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[16] ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_1_5), .B(\un1_add_reg_1_i[5] ), .C(
        I4_un1_CO1_i), .Y(\un3_addresult[5] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I14_S_0 (.A(\addresult_4[14] ), 
        .B(N254), .Y(\un3_addresult[14] ));
    OR2 \addresult_RNIQKFE[12]  (.A(\addresult_4[12] ), .B(N_254), .Y(
        N_91));
    OR2 \addresult_RNIF64E[6]  (.A(\addresult_4[6] ), .B(N_254), .Y(
        N_179));
    NOR3C un3_addresult_ADD_20x20_slow_I8_un1_CO1_0_m6 (.A(
        ADD_20x20_slow_I6_S_0_0), .B(ADD_20x20_slow_I8_un1_CO1_0_m6_0), 
        .C(ADD_20x20_slow_I7_S_0_0), .Y(
        ADD_20x20_slow_I8_un1_CO1_0_N_7_i));
    XOR2 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        ADD_20x20_slow_I4_S_0_0), .B(ADD_20x20_slow_I3_CO1_m12_0), .Y(
        \un3_addresult[4] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I18_S_0 (.A(\addresult_4[18] ), 
        .B(N270), .Y(\un3_addresult[18] ));
    AOI1B \addresult_RNIAA911[3]  (.A(\addresult_4[3] ), .B(N_273), .C(
        N_210_0), .Y(signal_data_iv_0_6_3));
    DFN1P0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .PRE(s_acq_change_0_s_rst), .Q(
        \un1_add_reg_1_i[5] ));
    AO1 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(\addresult_4[8] ), 
        .B(N240), .C(ADD_20x20_slow_I8_un1_CO1_0), .Y(I8_un1_CO1));
    NOR2A un3_addresult_ADD_20x20_slow_I1_un5_CO1_m2_0_a2_0 (.A(
        \addresult_4[0] ), .B(un1_n_s_change_0_1[0]), .Y(
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_0));
    OR2 \addresult_RNIII4E[9]  (.A(\addresult_4[9] ), .B(N_254), .Y(
        N_139));
    OAI1 un3_addresult_ADD_20x20_slow_I2_un1_CO1_0 (.A(N228), .B(
        un1_ten_choice_one_0_1_2), .C(\addresult_4[2] ), .Y(
        ADD_20x20_slow_I2_un1_CO1_0));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[2] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult_3[7] ), .C(un1_ten_choice_one_0_1_7), .Y(N240));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0_0 (.A(\addresult_4[6] ), 
        .B(un1_ten_choice_one_0_1_6), .Y(ADD_20x20_slow_I6_S_0_0));
    NOR2 un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_a5_2 (.A(N_216), .B(
        ADD_20x20_slow_I3_CO1tt_m1_0_a2), .Y(
        ADD_20x20_slow_I3_CO1_N_16));
    AO1A un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_0 (.A(
        \addresult_4[3] ), .B(un1_n_s_change_0_1[3]), .C(
        ADD_20x20_slow_I3_CO1_N_16), .Y(ADD_20x20_slow_I3_CO1_m12_0_0));
    OA1B un3_addresult_ADD_20x20_slow_I3_CO1tt_m1_0_a2 (.A(
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_2), .B(
        ADD_20x20_slow_I1_un3_CO1_m2_0_a2_2), .C(N_210), .Y(
        ADD_20x20_slow_I3_CO1tt_m1_0_a2));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e (.A(
        ADD_20x20_slow_I19_Y_0_m6_e_2), .B(
        ADD_20x20_slow_I19_Y_0_m6_e_1), .C(
        ADD_20x20_slow_I19_Y_0_m6_e_3), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_2_0));
    XNOR2 un3_addresult_ADD_20x20_slow_I16_S_0 (.A(\addresult_4[16] ), 
        .B(N262), .Y(\un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[3] ));
    OR2 \addresult_RNIPKFE[11]  (.A(\addresult_4[11] ), .B(N_254), .Y(
        N_155));
    NOR2A un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_o5 (.A(
        \addresult_4[3] ), .B(un1_n_s_change_0_1[3]), .Y(
        ADD_20x20_slow_I3_CO1_m12_0_o5));
    OA1 un3_addresult_ADD_20x20_slow_I9_CO1_0 (.A(I8_un1_CO1), .B(
        \addresult_4[9] ), .C(un1_ten_choice_one_0_1_9), .Y(
        ADD_20x20_slow_I9_CO1_0));
    AX1 un3_addresult_ADD_20x20_slow_I17_S_0 (.A(N262), .B(
        \addresult_4[16] ), .C(\addresult_4[17] ), .Y(
        \un3_addresult[17] ));
    OR2 \addresult_RNIHE4E[8]  (.A(\addresult_4[8] ), .B(N_254), .Y(
        N_131));
    OR3 \addresult_RNI4OGN[7]  (.A(\addresult_3[7] ), .B(
        \addresult_4[8] ), .C(un1_ten_choice_one_0_1_7), .Y(d_N_8_2));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[14] ));
    OA1B un3_addresult_ADD_20x20_slow_I1_CO1_0 (.A(
        ADD_20x20_slow_I1_un3_CO1_m2_0_a2_2), .B(
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_2), .C(N_210), .Y(
        ADD_20x20_slow_I1_CO1_0));
    AO1 un3_addresult_ADD_20x20_slow_I1_CO1 (.A(
        un1_ten_choice_one_0_1_1), .B(\addresult_4[1] ), .C(
        ADD_20x20_slow_I1_CO1_0), .Y(N228));
    XNOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(r_N_7_i), .B(
        \addresult_4[12] ), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    MX2C un3_addresult_ADD_20x20_slow_I8_un1_CO1_1 (.A(
        \addresult_RNIM85T1[7]_net_1 ), .B(r_N_2_1_i_0), .S(
        ADD_20x20_slow_I8_un1_CO1_0_N_7_i), .Y(
        ADD_20x20_slow_I8_un1_CO1_0));
    MIN3 un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(
        ADD_20x20_slow_I3_CO1_m12_0), .B(\addresult_4[4] ), .C(
        un1_ten_choice_one_0_1_4), .Y(I4_un1_CO1_i));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_1 (.A(
        \addresult_3[13] ), .B(\addresult_4[14] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_1));
    AO1 un3_addresult_ADD_20x20_slow_I10_un1_CO1_0_tz_0 (.A(
        \addresult_4[9] ), .B(I8_un1_CO1), .C(\addresult_4[10] ), .Y(
        ADD_20x20_slow_I10_un1_CO1_0_tz_0));
    AOI1B \addresult_RNI62911[1]  (.A(\addresult_4[1] ), .B(N_273), .C(
        N_243), .Y(signal_data_iv_0_0_6[1]));
    OR3 un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_a5_0_1 (.A(
        ADD_20x20_slow_I3_CO1_m3_e), .B(ADD_20x20_slow_I3_CO1_m12_0_o5)
        , .C(ADD_20x20_slow_I3_CO1_m12_0_o5_0), .Y(
        ADD_20x20_slow_I3_CO1_m12_0_a5_0_1));
    OR2 \addresult_RNITKFE[15]  (.A(\addresult_3[15] ), .B(N_254), .Y(
        N_115));
    NOR2A un3_addresult_ADD_20x20_slow_I3_CO1_m3_e (.A(
        \addresult_4[1] ), .B(un1_n_s_change_0_1[1]), .Y(
        ADD_20x20_slow_I3_CO1_m3_e));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_2 (.A(
        \addresult_3[15] ), .B(\addresult_4[16] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_2));
    OA1 un3_addresult_ADD_20x20_slow_I10_un1_CO1_0 (.A(
        ADD_20x20_slow_I9_CO1_0), .B(ADD_20x20_slow_I10_un1_CO1_0_tz_0)
        , .C(un1_ten_choice_one_0_1_10), .Y(
        ADD_20x20_slow_I10_un1_CO1_0));
    XOR2 un3_addresult_ADD_20x20_slow_I7_S_0_0 (.A(
        un1_ten_choice_one_0_1_7), .B(\addresult_3[7] ), .Y(
        ADD_20x20_slow_I7_S_0_0));
    OR3B un3_addresult_ADD_20x20_slow_I17_CO1 (.A(\addresult_4[16] ), 
        .B(\addresult_4[17] ), .C(N262), .Y(N270));
    NOR2A un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_o5_0 (.A(
        \addresult_4[2] ), .B(un1_n_s_change_0_1[2]), .Y(
        ADD_20x20_slow_I3_CO1_m12_0_o5_0));
    AX1 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(N254), .B(
        \addresult_4[14] ), .C(\addresult_3[15] ), .Y(
        \un3_addresult[15] ));
    OR2 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(I10_un5_CO1), .B(
        ADD_20x20_slow_I10_un1_CO1_0), .Y(I10_un1_CO1));
    NOR3B un3_addresult_ADD_20x20_slow_I1_un5_CO1_m2_0_a2_2 (.A(
        ADD_20x20_slow_I1_un5_CO1_m2_0_a2_0), .B(\addresult_4[1] ), .C(
        N_213), .Y(ADD_20x20_slow_I1_un5_CO1_m2_0_a2_2));
    OR3A \addresult_RNIIUVI[16]  (.A(\addresult_4[16] ), .B(N_249_0), 
        .C(N_251), .Y(N_192));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[11] ));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[17] ));
    AO1 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(\addresult_4[9] ), .B(
        I8_un1_CO1), .C(ADD_20x20_slow_I9_CO1_0), .Y(N244));
    NOR2B un3_addresult_ADD_20x20_slow_I10_un5_CO1 (.A(
        \addresult_4[10] ), .B(N244), .Y(I10_un5_CO1));
    OR2A \addresult_RNIE24E[5]  (.A(\un1_add_reg_1_i[5] ), .B(N_254), 
        .Y(N_171));
    AOI1B \addresult_RNI86911[2]  (.A(\addresult_4[2] ), .B(N_273), .C(
        N_226), .Y(signal_data_iv_0_6_2));
    MAJ3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult_4[6] ), .C(un1_ten_choice_one_0_1_6), .Y(I6_un1_CO1)
        );
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_1_10), .B(\addresult_4[10] ), .C(N244), 
        .Y(\un3_addresult[10] ));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[7] ));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_3 (.A(
        \addresult_4[12] ), .B(\addresult_4[18] ), .C(
        \addresult_4[17] ), .Y(ADD_20x20_slow_I19_Y_0_m6_e_3));
    AX1 un3_addresult_ADD_20x20_slow_I13_S_0 (.A(r_N_7_i), .B(
        \addresult_4[12] ), .C(\addresult_3[13] ), .Y(
        \un3_addresult[13] ));
    OR3C \addresult_RNIM85T1[7]  (.A(d_N_8_2), .B(
        un1_ten_choice_one_0_1_8), .C(d_N_7_2), .Y(
        \addresult_RNIM85T1[7]_net_1 ));
    MAJ3 \addresult_RNI0GEU5[5]  (.A(I4_un1_CO1_i), .B(
        \un1_add_reg_1_i[5] ), .C(un1_ten_choice_one_0_1_5), .Y(
        r_N_2_1_i_0));
    AX1C un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        ADD_20x20_slow_I2_un1_CO1_0), .B(I2_un4_CO1), .C(
        ADD_20x20_slow_I3_S_0_0), .Y(\un3_addresult[3] ));
    NOR3A un3_addresult_ADD_20x20_slow_I3_CO1_m12_0_a5 (.A(
        un1_n_s_change_0_1[2]), .B(\addresult_4[2] ), .C(
        ADD_20x20_slow_I3_CO1_N_9), .Y(ADD_20x20_slow_I3_CO1_m12_0_a5));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[18] ));
    OR3A \addresult_RNIKUVI[18]  (.A(\addresult_4[18] ), .B(N_249), .C(
        N_251), .Y(N_224));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        ADD_20x20_slow_I6_S_0_0), .B(N236), .Y(\un3_addresult[6] ));
    OR3A \addresult_RNIJUVI[17]  (.A(\addresult_4[17] ), .B(N_249_0), 
        .C(N_251), .Y(N_241));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[13] ));
    XOR2 un3_addresult_ADD_20x20_slow_I1_S_0_0 (.A(\addresult_4[1] ), 
        .B(un1_ten_choice_one_0_1_1), .Y(ADD_20x20_slow_I1_S_0_0));
    OR3A \addresult_RNILUVI[19]  (.A(\addresult_4[19] ), .B(N_249_0), 
        .C(N_251), .Y(N_208));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[9] ));
    DFN1E1C0 \addresult[19]  (.D(\addresult_RNO_2[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .E(
        ADD_20x20_slow_I19_Y_0_m6_e_2_0), .Q(\addresult_4[19] ));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[0] ));
    NOR2A un3_addresult_ADD_20x20_slow_I8_un1_CO1_0_m6_0 (.A(
        un1_ten_choice_one_0_1_8), .B(\addresult_4[8] ), .Y(
        ADD_20x20_slow_I8_un1_CO1_0_m6_0));
    XOR2 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(I6_un1_CO1), .B(
        ADD_20x20_slow_I7_S_0_0), .Y(\un3_addresult[7] ));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_1_9), .B(\addresult_4[9] ), .C(I8_un1_CO1)
        , .Y(\un3_addresult[9] ));
    XOR3 un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        un1_ten_choice_one_0_1_2), .B(\addresult_4[2] ), .C(N228), .Y(
        \un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    XOR2 un3_addresult_ADD_20x20_slow_I11_S_0_0 (.A(\addresult_4[11] ), 
        .B(un1_ten_choice_one_0_1_11), .Y(ADD_20x20_slow_I11_S_0_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_4[1] ));
    
endmodule


module add_reg_add_reg_2_6(
       addresult_RNIJE5C,
       addresult_RNIFE5C,
       addresult_RNIBOIB,
       addresult_0_15,
       addresult_0_13,
       signal_data_iv_0_0_1,
       signal_data_iv_0_1_0,
       signal_data_iv_0_1_3,
       signal_data_iv_0_1_2,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_6,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_214,
       N_182,
       N_221,
       N_249,
       N_198,
       N_256,
       N_249_0,
       N_231,
       N_174,
       N_158,
       N_150,
       N_134,
       N_126,
       N_118,
       N_255,
       N_86,
       N_210,
       N_212,
       N_184,
       N_233,
       N_200,
       N_216,
       N_270
    );
output [14:14] addresult_RNIJE5C;
output [10:10] addresult_RNIFE5C;
output [5:5] addresult_RNIBOIB;
output addresult_0_15;
output addresult_0_13;
output [1:1] signal_data_iv_0_0_1;
output signal_data_iv_0_1_0;
output signal_data_iv_0_1_3;
output signal_data_iv_0_1_2;
input  [2:0] un1_n_s_change_0_1;
input  [11:1] un1_ten_choice_one_0_6;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
output N_214;
output N_182;
input  N_221;
input  N_249;
output N_198;
input  N_256;
input  N_249_0;
output N_231;
output N_174;
output N_158;
output N_150;
output N_134;
output N_126;
output N_118;
input  N_255;
output N_86;
input  N_210;
input  N_212;
input  N_184;
input  N_233;
input  N_200;
input  N_216;
input  N_270;

    wire ADD_20x20_slow_I7_CO1_0_tz_0, \addresult_0[6] , N236, 
        \addresult_0[7] , ADD_20x20_slow_I6_S_0_0, 
        ADD_20x20_slow_I5_CO1_0_tz_0, I4_un5_CO1, \addresult_0[5] , 
        ADD_20x20_slow_I2_un1_CO1_m4_i_0, ADD_20x20_slow_I1_CO1_m5_i_0, 
        \addresult_0[2] , \addresult_0[3] , \addresult_0[1] , 
        \addresult_0[0] , \un3_addresult[11] , \addresult_0[11] , 
        I10_un1_CO1, \un3_addresult[9] , \addresult_0[9] , I8_un1_CO1, 
        \un3_addresult[8] , \addresult_0[8] , N240, \un3_addresult[7] , 
        I6_un1_CO1, \un3_addresult[6] , \un3_addresult[5] , I4_un1_CO1, 
        \un3_addresult[4] , \addresult_0[4] , N232, \un3_addresult[3] , 
        ADD_20x20_slow_I2_un1_CO1_N_5, \un3_addresult[10] , 
        \addresult_0[10] , N244, \un3_addresult[1] , I0_un1_CO1, 
        \un3_addresult[2] , ADD_20x20_slow_I1_CO1_m5_i_0_0, 
        ADD_20x20_slow_I7_CO1_0_tz, ADD_20x20_slow_I6_un1_CO1_0, 
        ADD_20x20_slow_I1_CO1tt_m1_e_0, ADD_20x20_slow_I5_CO1_0, 
        ADD_20x20_slow_I4_un1_CO1_0, I5_un5_CO1, I7_un5_CO1, N248, 
        N254, \addresult_0[12] , \un3_addresult[12] , 
        \un3_addresult[13] , \un3_addresult[14] , \addresult_0[14] , 
        \un3_addresult[18] , \addresult_0[18] , N270, 
        \un3_addresult[19] , \addresult_0[19] , \un3_addresult[17] , 
        N262, \addresult_0[16] , \addresult_0[17] , 
        \un3_addresult[15] , \un3_addresult[0] , \un3_addresult[16] , 
        GND, VCC, GND_0, VCC_0;
    
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        un1_ten_choice_one_0_6[11]), .B(\addresult_0[11] ), .C(
        I10_un1_CO1), .Y(\un3_addresult[11] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[12] ));
    AO1 un3_addresult_ADD_20x20_slow_I7_CO1_0_tz_0 (.A(
        \addresult_0[6] ), .B(N236), .C(\addresult_0[7] ), .Y(
        ADD_20x20_slow_I7_CO1_0_tz_0));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_6[8]), .B(\addresult_0[8] ), .C(N240), .Y(
        \un3_addresult[8] ));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[10] ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[6] ));
    AO13 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(
        un1_ten_choice_one_0_6[3]), .B(\addresult_0[3] ), .C(
        ADD_20x20_slow_I2_un1_CO1_N_5), .Y(N232));
    AOI1B \addresult_RNIODDS[0]  (.A(\addresult_0[0] ), .B(N_270), .C(
        N_184), .Y(signal_data_iv_0_1_0));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[8] ));
    NOR2A un3_addresult_ADD_20x20_slow_I1_CO1tt_m1_e (.A(
        \addresult_0[0] ), .B(un1_n_s_change_0_1[0]), .Y(
        ADD_20x20_slow_I1_CO1tt_m1_e_0));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(I0_un1_CO1), .B(
        \addresult_0[1] ), .C(un1_ten_choice_one_0_6[1]), .Y(
        \un3_addresult[1] ));
    OR2 \addresult_RNIGE5C[11]  (.A(\addresult_0[11] ), .B(N_255), .Y(
        N_150));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_0_15));
    OR2 \addresult_RNID0JB[7]  (.A(\addresult_0[7] ), .B(N_255), .Y(
        N_118));
    VCC VCC_i (.Y(VCC));
    AO1B un3_addresult_ADD_20x20_slow_I5_CO1_0 (.A(
        ADD_20x20_slow_I5_CO1_0_tz_0), .B(ADD_20x20_slow_I4_un1_CO1_0), 
        .C(un1_ten_choice_one_0_6[5]), .Y(ADD_20x20_slow_I5_CO1_0));
    MAJ3 un3_addresult_ADD_20x20_slow_I11_CO1 (.A(I10_un1_CO1), .B(
        \addresult_0[11] ), .C(un1_ten_choice_one_0_6[11]), .Y(N248));
    OR2B un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I5_un5_CO1), .B(
        ADD_20x20_slow_I5_CO1_0), .Y(N236));
    OA1 un3_addresult_ADD_20x20_slow_I6_un1_CO1_0 (.A(N236), .B(
        \addresult_0[6] ), .C(un1_ten_choice_one_0_6[6]), .Y(
        ADD_20x20_slow_I6_un1_CO1_0));
    OR2 \addresult_RNIJE5C[14]  (.A(\addresult_0[14] ), .B(N_255), .Y(
        addresult_RNIJE5C[14]));
    OR3A \addresult_RNIBOLG[18]  (.A(\addresult_0[18] ), .B(N_249), .C(
        N_256), .Y(N_214));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[4] ));
    NOR3B un3_addresult_ADD_20x20_slow_I15_CO1 (.A(\addresult_0[14] ), 
        .B(addresult_0_15), .C(N254), .Y(N262));
    AX1B un3_addresult_ADD_20x20_slow_I0_S_0 (.A(N_221), .B(
        un1_n_s_change_0_1[0]), .C(\addresult_0[0] ), .Y(
        \un3_addresult[0] ));
    OR3C un3_addresult_ADD_20x20_slow_I13_CO1 (.A(N248), .B(
        \addresult_0[12] ), .C(addresult_0_13), .Y(N254));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[16] ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_6[5]), .B(\addresult_0[5] ), .C(
        I4_un1_CO1), .Y(\un3_addresult[5] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I14_S_0 (.A(\addresult_0[14] ), 
        .B(N254), .Y(\un3_addresult[14] ));
    XOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0_6[4]), .B(\addresult_0[4] ), .C(N232), .Y(
        \un3_addresult[4] ));
    XOR2 un3_addresult_ADD_20x20_slow_I18_S_0 (.A(\addresult_0[18] ), 
        .B(N270), .Y(\un3_addresult[18] ));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[5] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_0[8] ), .C(un1_ten_choice_one_0_6[8]), .Y(
        I8_un1_CO1));
    OR2 un3_addresult_ADD_20x20_slow_I7_CO1_0_tz (.A(
        ADD_20x20_slow_I7_CO1_0_tz_0), .B(ADD_20x20_slow_I6_un1_CO1_0), 
        .Y(ADD_20x20_slow_I7_CO1_0_tz));
    AX1C un3_addresult_ADD_20x20_slow_I19_Y_0 (.A(N270), .B(
        \addresult_0[18] ), .C(\addresult_0[19] ), .Y(
        \un3_addresult[19] ));
    AO13 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m4_i_0 (.A(
        ADD_20x20_slow_I1_CO1_m5_i_0), .B(\addresult_0[2] ), .C(
        un1_n_s_change_0_1[2]), .Y(ADD_20x20_slow_I2_un1_CO1_m4_i_0));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[2] ));
    AO1B un3_addresult_ADD_20x20_slow_I7_CO1 (.A(
        un1_ten_choice_one_0_6[7]), .B(ADD_20x20_slow_I7_CO1_0_tz), .C(
        I7_un5_CO1), .Y(N240));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0_0 (.A(\addresult_0[6] ), 
        .B(un1_ten_choice_one_0_6[6]), .Y(ADD_20x20_slow_I6_S_0_0));
    OR2 \addresult_RNIFE5C[10]  (.A(\addresult_0[10] ), .B(N_255), .Y(
        addresult_RNIFE5C[10]));
    OR3A \addresult_RNICOLG[19]  (.A(\addresult_0[19] ), .B(N_249), .C(
        N_256), .Y(N_198));
    OR2B un3_addresult_ADD_20x20_slow_I5_un5_CO1 (.A(\addresult_0[5] ), 
        .B(I4_un1_CO1), .Y(I5_un5_CO1));
    XOR2 un3_addresult_ADD_20x20_slow_I16_S_0 (.A(\addresult_0[16] ), 
        .B(N262), .Y(\un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[3] ));
    AOI1B \addresult_RNIQHDS[1]  (.A(\addresult_0[1] ), .B(N_270), .C(
        N_233), .Y(signal_data_iv_0_0_1[1]));
    AOI1B \addresult_RNIUPDS[3]  (.A(\addresult_0[3] ), .B(N_270), .C(
        N_200), .Y(signal_data_iv_0_1_3));
    AX1C un3_addresult_ADD_20x20_slow_I17_S_0 (.A(N262), .B(
        \addresult_0[16] ), .C(\addresult_0[17] ), .Y(
        \un3_addresult[17] ));
    OR3A \addresult_RNIAOLG[17]  (.A(\addresult_0[17] ), .B(N_249_0), 
        .C(N_256), .Y(N_231));
    OR3A un3_addresult_ADD_20x20_slow_I1_CO1_m5_i (.A(
        ADD_20x20_slow_I1_CO1_m5_i_0), .B(N_212), .C(N_210), .Y(
        ADD_20x20_slow_I1_CO1_m5_i_0_0));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[14] ));
    XOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(\addresult_0[12] ), 
        .B(N248), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    OR3A \addresult_RNI9OLG[16]  (.A(\addresult_0[16] ), .B(N_249), .C(
        N_256), .Y(N_182));
    OR2 \addresult_RNICSIB[6]  (.A(\addresult_0[6] ), .B(N_255), .Y(
        N_174));
    OR2 \addresult_RNIAKIB[4]  (.A(\addresult_0[4] ), .B(N_255), .Y(
        N_158));
    OR2B un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(I4_un5_CO1), .B(
        ADD_20x20_slow_I4_un1_CO1_0), .Y(I4_un1_CO1));
    AOI1B \addresult_RNISLDS[2]  (.A(\addresult_0[2] ), .B(N_270), .C(
        N_216), .Y(signal_data_iv_0_1_2));
    NOR3C un3_addresult_ADD_20x20_slow_I17_CO1 (.A(N262), .B(
        \addresult_0[16] ), .C(\addresult_0[17] ), .Y(N270));
    OR2 \addresult_RNIBOIB[5]  (.A(\addresult_0[5] ), .B(N_255), .Y(
        addresult_RNIBOIB[5]));
    AX1 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(N254), .B(
        \addresult_0[14] ), .C(addresult_0_15), .Y(\un3_addresult[15] )
        );
    OR3A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m4_i (.A(
        ADD_20x20_slow_I2_un1_CO1_m4_i_0), .B(N_212), .C(N_210), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_5));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult_0[10] ), .C(un1_ten_choice_one_0_6[10]), .Y(
        I10_un1_CO1));
    OR2 \addresult_RNIE4JB[8]  (.A(\addresult_0[8] ), .B(N_255), .Y(
        N_126));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[11] ));
    OAI1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0 (.A(N232), .B(
        \addresult_0[4] ), .C(un1_ten_choice_one_0_6[4]), .Y(
        ADD_20x20_slow_I4_un1_CO1_0));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[17] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1), .B(
        \addresult_0[9] ), .C(un1_ten_choice_one_0_6[9]), .Y(N244));
    OR2 \addresult_RNIF8JB[9]  (.A(\addresult_0[9] ), .B(N_255), .Y(
        N_134));
    NOR2A un3_addresult_ADD_20x20_slow_I5_CO1_0_tz_0 (.A(I4_un5_CO1), 
        .B(\addresult_0[5] ), .Y(ADD_20x20_slow_I5_CO1_0_tz_0));
    OR2 \addresult_RNIHE5C[12]  (.A(\addresult_0[12] ), .B(N_255), .Y(
        N_86));
    AO1 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(\addresult_0[6] ), 
        .B(N236), .C(ADD_20x20_slow_I6_un1_CO1_0), .Y(I6_un1_CO1));
    OR2B un3_addresult_ADD_20x20_slow_I4_un5_CO1 (.A(\addresult_0[4] ), 
        .B(N232), .Y(I4_un5_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_6[10]), .B(\addresult_0[10] ), .C(N244), 
        .Y(\un3_addresult[10] ));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[7] ));
    OR2B un3_addresult_ADD_20x20_slow_I7_un5_CO1 (.A(\addresult_0[7] ), 
        .B(I6_un1_CO1), .Y(I7_un5_CO1));
    AX1C un3_addresult_ADD_20x20_slow_I13_S_0 (.A(N248), .B(
        \addresult_0[12] ), .C(addresult_0_13), .Y(\un3_addresult[13] )
        );
    XNOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        ADD_20x20_slow_I2_un1_CO1_N_5), .B(\addresult_0[3] ), .C(
        un1_ten_choice_one_0_6[3]), .Y(\un3_addresult[3] ));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[18] ));
    XOR2 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        ADD_20x20_slow_I6_S_0_0), .B(N236), .Y(\un3_addresult[6] ));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_0_13));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[9] ));
    DFN1C0 \addresult[19]  (.D(\un3_addresult[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[19] ));
    AO13 un3_addresult_ADD_20x20_slow_I1_CO1_m5_i_0 (.A(
        ADD_20x20_slow_I1_CO1tt_m1_e_0), .B(\addresult_0[1] ), .C(
        un1_n_s_change_0_1[1]), .Y(ADD_20x20_slow_I1_CO1_m5_i_0));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[0] ));
    OR3A un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(\addresult_0[0] ), 
        .B(N_221), .C(un1_n_s_change_0_1[0]), .Y(I0_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0_6[7]), .B(\addresult_0[7] ), .C(
        I6_un1_CO1), .Y(\un3_addresult[7] ));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_6[9]), .B(\addresult_0[9] ), .C(
        I8_un1_CO1), .Y(\un3_addresult[9] ));
    XOR3 un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        ADD_20x20_slow_I1_CO1_m5_i_0_0), .B(\addresult_0[2] ), .C(
        un1_ten_choice_one_0_6[2]), .Y(\un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_0[1] ));
    
endmodule


module add_reg_add_reg_2_5(
       s_addchoice,
       signal_data_iv_0_0_13,
       signal_data_en,
       signal_data_iv_0_13_2,
       signal_data_iv_0_13_3,
       signal_data_iv_0_13_0,
       un1_signal_acq_0,
       dataeight_0_a2_0_0,
       signal_data_0_iv_i_0,
       signal_data_iv_0_0_9,
       signal_data_iv_0_0_1,
       signal_data_iv_0_9_0,
       signal_data_iv_0_9_3,
       signal_data_iv_0_9_2,
       signal_data_iv_0_1_0,
       signal_data_iv_0_1_3,
       signal_data_iv_0_1_2,
       addresult_14,
       addresult_13,
       addresult_15,
       addresult_12,
       un1_ten_choice_one_0_7_2,
       un1_ten_choice_one_0_7_3,
       un1_ten_choice_one_0_7_5,
       un1_ten_choice_one_0_7_6,
       un1_ten_choice_one_0_7_7,
       un1_ten_choice_one_0_7_8,
       un1_ten_choice_one_0_7_9,
       un1_ten_choice_one_0_7_10,
       un1_ten_choice_one_0_7_11,
       un1_ten_choice_one_0_7_0,
       un1_n_s_change_0_1,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_228,
       N_245,
       N_196,
       G_1_0_a2_0,
       N_212,
       N_213,
       N_182,
       N_33,
       N_256,
       N_231,
       N_198,
       N_214,
       N_267,
       N_220
    );
input  [0:0] s_addchoice;
input  [1:1] signal_data_iv_0_0_13;
input  [9:9] signal_data_en;
input  signal_data_iv_0_13_2;
input  signal_data_iv_0_13_3;
input  signal_data_iv_0_13_0;
output [3:0] un1_signal_acq_0;
input  [0:0] dataeight_0_a2_0_0;
output [11:4] signal_data_0_iv_i_0;
input  [1:1] signal_data_iv_0_0_9;
input  [1:1] signal_data_iv_0_0_1;
input  signal_data_iv_0_9_0;
input  signal_data_iv_0_9_3;
input  signal_data_iv_0_9_2;
input  signal_data_iv_0_1_0;
input  signal_data_iv_0_1_3;
input  signal_data_iv_0_1_2;
output addresult_14;
output addresult_13;
output addresult_15;
output addresult_12;
input  un1_ten_choice_one_0_7_2;
input  un1_ten_choice_one_0_7_3;
input  un1_ten_choice_one_0_7_5;
input  un1_ten_choice_one_0_7_6;
input  un1_ten_choice_one_0_7_7;
input  un1_ten_choice_one_0_7_8;
input  un1_ten_choice_one_0_7_9;
input  un1_ten_choice_one_0_7_10;
input  un1_ten_choice_one_0_7_11;
input  un1_ten_choice_one_0_7_0;
input  [4:0] un1_n_s_change_0_1;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
output N_228;
output N_245;
output N_196;
input  G_1_0_a2_0;
output N_212;
input  N_213;
input  N_182;
input  N_33;
input  N_256;
input  N_231;
input  N_198;
input  N_214;
input  N_267;
input  N_220;

    wire ADD_20x20_slow_I4_S_0_0, \addresult[4]_net_1 , 
        ADD_20x20_slow_I4_un1_CO1_m11_i_0, \addresult[2]_net_1 , 
        ADD_20x20_slow_I1_S_0_0, \addresult[0]_net_1 , 
        \addresult[1]_net_1 , ADD_20x20_slow_I1_CO1_m5_i_0, 
        ADD_20x20_slow_I1_CO1tt_m1_e, ADD_20x20_slow_I19_Y_0_m6_e_3, 
        \addresult[18]_net_1 , \addresult[17]_net_1 , 
        ADD_20x20_slow_I19_Y_0_m6_e_2, \addresult[16]_net_1 , 
        ADD_20x20_slow_I19_Y_0_m6_e_1, \signal_data_iv_0_12[2] , 
        \signal_data_iv_0_0[2] , \signal_data_iv_0_12[3] , 
        \signal_data_iv_0_0[3] , \addresult[3]_net_1 , 
        \signal_data_iv_0_0_12[1] , \signal_data_iv_0_0_0[1] , 
        \addresult[5]_net_1 , \addresult[11]_net_1 , 
        \addresult[7]_net_1 , \addresult[8]_net_1 , 
        \addresult[9]_net_1 , \addresult[10]_net_1 , 
        \addresult[6]_net_1 , \signal_data_iv_0_12[0] , 
        \signal_data_iv_0_0[0] , ADD_20x20_slow_I19_Y_0_m6_e, 
        \un3_addresult[11] , I10_un1_CO1, \un3_addresult[10] , N244, 
        \un3_addresult[9] , I8_un1_CO1, \un3_addresult[8] , N240, 
        \un3_addresult[7] , I6_un1_CO1, \un3_addresult[6] , N236, 
        \un3_addresult[5] , I4_un1_CO1, \un3_addresult[4] , N232, 
        \un3_addresult[3] , I2_un1_CO1, \un3_addresult[1] , 
        \un3_addresult[2] , ADD_20x20_slow_I1_CO1_m5_i, 
        ADD_20x20_slow_I4_un1_CO1_m11_i, 
        ADD_20x20_slow_I4_un1_CO1_N_14_i_i, 
        ADD_20x20_slow_I4_un1_CO1_N_15_i_i, 
        ADD_20x20_slow_I2_un1_CO1_0_tz, \addresult_RNO[19]_net_1 , 
        r_N_7_2_i, \addresult[19]_net_1 , I2_un3_CO1_i, 
        \addresult_RNIUESN[4]_net_1 , d_N_13, d_N_4, N254, 
        \un3_addresult[12] , \un3_addresult[13] , \un3_addresult[14] , 
        \un3_addresult[0] , \un3_addresult[15] , N262, I16_un1_CO1, 
        \un3_addresult[16] , \un3_addresult[17] , \un3_addresult[18] , 
        GND, VCC, GND_0, VCC_0;
    
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        un1_ten_choice_one_0_7_11), .B(\addresult[11]_net_1 ), .C(
        I10_un1_CO1), .Y(\un3_addresult[11] ));
    OR3B \addresult_RNIKG0D[16]  (.A(G_1_0_a2_0), .B(
        \addresult[16]_net_1 ), .C(s_addchoice[0]), .Y(N_196));
    AOI1B \addresult_RNI0P1T[2]  (.A(\addresult[2]_net_1 ), .B(N_267), 
        .C(N_214), .Y(\signal_data_iv_0_0[2] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_12));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_7_8), .B(\addresult[8]_net_1 ), .C(N240), 
        .Y(\un3_addresult[8] ));
    AOI1 \addresult_RNIQAPS7[1]  (.A(signal_data_iv_0_0_13[1]), .B(
        \signal_data_iv_0_0_12[1] ), .C(signal_data_en[9]), .Y(
        un1_signal_acq_0[1]));
    NOR3C \addresult_RNI01EG3[1]  (.A(signal_data_iv_0_0_1[1]), .B(
        \signal_data_iv_0_0_0[1] ), .C(signal_data_iv_0_0_9[1]), .Y(
        \signal_data_iv_0_0_12[1] ));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[10]_net_1 ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[6]_net_1 ));
    AX1B un3_addresult_ADD_20x20_slow_I4_un1_CO1_m11_i_x2_0 (.A(N_220), 
        .B(un1_n_s_change_0_1[3]), .C(\addresult[3]_net_1 ), .Y(
        ADD_20x20_slow_I4_un1_CO1_N_15_i_i));
    MAJ3 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(I2_un1_CO1), .B(
        \addresult[3]_net_1 ), .C(un1_ten_choice_one_0_7_3), .Y(N232));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[8]_net_1 ));
    NOR2A un3_addresult_ADD_20x20_slow_I1_CO1tt_m1_e (.A(
        \addresult[0]_net_1 ), .B(un1_n_s_change_0_1[0]), .Y(
        ADD_20x20_slow_I1_CO1tt_m1_e));
    AX1D un3_addresult_ADD_20x20_slow_I4_S_0_0 (.A(N_220), .B(
        un1_n_s_change_0_1[4]), .C(\addresult[4]_net_1 ), .Y(
        ADD_20x20_slow_I4_S_0_0));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1_0_tz (.A(
        un1_n_s_change_0_1[2]), .B(\addresult[2]_net_1 ), .Y(
        ADD_20x20_slow_I2_un1_CO1_0_tz));
    AX1D un3_addresult_ADD_20x20_slow_I1_S_0 (.A(N_220), .B(
        un1_n_s_change_0_1[1]), .C(ADD_20x20_slow_I1_S_0_0), .Y(
        \un3_addresult[1] ));
    OA1B \addresult_RNIROCC[8]  (.A(N_256), .B(\addresult[8]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[8]));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_15));
    OR2A un3_addresult_ADD_20x20_slow_I2_un3_CO1 (.A(
        \addresult[2]_net_1 ), .B(un1_ten_choice_one_0_7_2), .Y(
        I2_un3_CO1_i));
    XNOR2 \addresult_RNO[19]  (.A(r_N_7_2_i), .B(\addresult[19]_net_1 )
        , .Y(\addresult_RNO[19]_net_1 ));
    OAI1 un3_addresult_ADD_20x20_slow_I2_un1_CO1 (.A(
        ADD_20x20_slow_I1_CO1_m5_i), .B(ADD_20x20_slow_I2_un1_CO1_0_tz)
        , .C(I2_un3_CO1_i), .Y(I2_un1_CO1));
    VCC VCC_i (.Y(VCC));
    MAJ3 un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I4_un1_CO1), .B(
        \addresult[5]_net_1 ), .C(un1_ten_choice_one_0_7_5), .Y(N236));
    OA1B \addresult_RNIEG0D[10]  (.A(N_256), .B(\addresult[10]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[10]));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[4]_net_1 ));
    AX1B un3_addresult_ADD_20x20_slow_I4_un1_CO1_m11_i_x2 (.A(N_220), 
        .B(un1_n_s_change_0_1[4]), .C(\addresult[4]_net_1 ), .Y(
        ADD_20x20_slow_I4_un1_CO1_N_14_i_i));
    OR3B un3_addresult_ADD_20x20_slow_I15_CO1 (.A(addresult_14), .B(
        addresult_15), .C(N254), .Y(N262));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0_7_0), .B(\addresult[0]_net_1 ), .Y(
        \un3_addresult[0] ));
    OR3B un3_addresult_ADD_20x20_slow_I13_CO1 (.A(addresult_12), .B(
        addresult_13), .C(r_N_7_2_i), .Y(N254));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[16]_net_1 ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_7_5), .B(\addresult[5]_net_1 ), .C(
        I4_un1_CO1), .Y(\un3_addresult[5] ));
    XNOR2 un3_addresult_ADD_20x20_slow_I14_S_0 (.A(addresult_14), .B(
        N254), .Y(\un3_addresult[14] ));
    OR3B \addresult_RNILG0D[17]  (.A(G_1_0_a2_0), .B(
        \addresult[17]_net_1 ), .C(s_addchoice[0]), .Y(N_245));
    NOR3C \addresult_RNIG1FG3[3]  (.A(signal_data_iv_0_1_3), .B(
        \signal_data_iv_0_0[3] ), .C(signal_data_iv_0_9_3), .Y(
        \signal_data_iv_0_12[3] ));
    AOI1 \addresult_RNIAAOS7[0]  (.A(signal_data_iv_0_13_0), .B(
        \signal_data_iv_0_12[0] ), .C(signal_data_en[9]), .Y(
        un1_signal_acq_0[0]));
    XNOR2 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        ADD_20x20_slow_I4_S_0_0), .B(N232), .Y(\un3_addresult[4] ));
    AX1C un3_addresult_ADD_20x20_slow_I18_S_0 (.A(I16_un1_CO1), .B(
        \addresult[17]_net_1 ), .C(\addresult[18]_net_1 ), .Y(
        \un3_addresult[18] ));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[5]_net_1 ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult[8]_net_1 ), .C(un1_ten_choice_one_0_7_8), .Y(
        I8_un1_CO1));
    NOR3C \addresult_RNIOGDG3[0]  (.A(signal_data_iv_0_1_0), .B(
        \signal_data_iv_0_0[0] ), .C(signal_data_iv_0_9_0), .Y(
        \signal_data_iv_0_12[0] ));
    OR3B \addresult_RNIMG0D[18]  (.A(G_1_0_a2_0), .B(
        \addresult[18]_net_1 ), .C(s_addchoice[0]), .Y(N_228));
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[2]_net_1 ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult[7]_net_1 ), .C(un1_ten_choice_one_0_7_7), .Y(N240));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e (.A(
        ADD_20x20_slow_I19_Y_0_m6_e_2), .B(
        ADD_20x20_slow_I19_Y_0_m6_e_1), .C(
        ADD_20x20_slow_I19_Y_0_m6_e_3), .Y(ADD_20x20_slow_I19_Y_0_m6_e)
        );
    OA1B \addresult_RNIN8CC[4]  (.A(N_256), .B(\addresult[4]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[4]));
    XNOR2 un3_addresult_ADD_20x20_slow_I16_S_0 (.A(
        \addresult[16]_net_1 ), .B(N262), .Y(\un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[3]_net_1 ));
    AOI1B \addresult_RNISG1T[0]  (.A(\addresult[0]_net_1 ), .B(N_267), 
        .C(N_182), .Y(\signal_data_iv_0_0[0] ));
    XOR2 un3_addresult_ADD_20x20_slow_I17_S_0 (.A(
        \addresult[17]_net_1 ), .B(I16_un1_CO1), .Y(
        \un3_addresult[17] ));
    OR3 un3_addresult_ADD_20x20_slow_I1_CO1_m5_i (.A(
        dataeight_0_a2_0_0[0]), .B(ADD_20x20_slow_I1_CO1_m5_i_0), .C(
        N_213), .Y(ADD_20x20_slow_I1_CO1_m5_i));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_14));
    XNOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(r_N_7_2_i), .B(
        addresult_12), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_1 (.A(addresult_13)
        , .B(addresult_14), .Y(ADD_20x20_slow_I19_Y_0_m6_e_1));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_2 (.A(addresult_15)
        , .B(\addresult[16]_net_1 ), .Y(ADD_20x20_slow_I19_Y_0_m6_e_2));
    NOR2A un3_addresult_ADD_20x20_slow_I16_un1_CO1 (.A(
        \addresult[16]_net_1 ), .B(N262), .Y(I16_un1_CO1));
    AX1 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(N254), .B(
        addresult_14), .C(addresult_15), .Y(\un3_addresult[15] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult[10]_net_1 ), .C(un1_ten_choice_one_0_7_10), .Y(
        I10_un1_CO1));
    OR2A \addresult_RNIUESN[4]  (.A(d_N_13), .B(N_220), .Y(
        \addresult_RNIUESN[4]_net_1 ));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[11]_net_1 ));
    OR3C un3_addresult_ADD_20x20_slow_I4_un1_CO1_m11_i (.A(
        ADD_20x20_slow_I4_un1_CO1_N_14_i_i), .B(
        ADD_20x20_slow_I4_un1_CO1_m11_i_0), .C(
        ADD_20x20_slow_I4_un1_CO1_N_15_i_i), .Y(
        ADD_20x20_slow_I4_un1_CO1_m11_i));
    AOI1B \addresult_RNIUK1T[1]  (.A(\addresult[1]_net_1 ), .B(N_267), 
        .C(N_231), .Y(\signal_data_iv_0_0_0[1] ));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[17]_net_1 ));
    MAJ3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1), .B(
        \addresult[9]_net_1 ), .C(un1_ten_choice_one_0_7_9), .Y(N244));
    OA1B \addresult_RNIPGCC[6]  (.A(N_256), .B(\addresult[6]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[6]));
    AOI1B \addresult_RNI2T1T[3]  (.A(\addresult[3]_net_1 ), .B(N_267), 
        .C(N_198), .Y(\signal_data_iv_0_0[3] ));
    AXO6 un3_addresult_ADD_20x20_slow_I4_un1_CO1_m11_i_0 (.A(N_220), 
        .B(un1_n_s_change_0_1[2]), .C(\addresult[2]_net_1 ), .Y(
        ADD_20x20_slow_I4_un1_CO1_m11_i_0));
    AOI1 \addresult_RNIABQS7[2]  (.A(signal_data_iv_0_13_2), .B(
        \signal_data_iv_0_12[2] ), .C(signal_data_en[9]), .Y(
        un1_signal_acq_0[2]));
    OA1B \addresult_RNIFG0D[11]  (.A(N_256), .B(\addresult[11]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[11]));
    AO13 \addresult_RNIDE0E[3]  (.A(un1_n_s_change_0_1[3]), .B(
        un1_n_s_change_0_1[2]), .C(\addresult[3]_net_1 ), .Y(d_N_4));
    MAJ3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult[6]_net_1 ), .C(un1_ten_choice_one_0_7_6), .Y(
        I6_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_7_10), .B(\addresult[10]_net_1 ), .C(N244)
        , .Y(\un3_addresult[10] ));
    OA1B \addresult_RNIOCCC[5]  (.A(N_256), .B(\addresult[5]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[5]));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[7]_net_1 ));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_3 (.A(addresult_12)
        , .B(\addresult[18]_net_1 ), .C(\addresult[17]_net_1 ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_3));
    AX1 un3_addresult_ADD_20x20_slow_I13_S_0 (.A(r_N_7_2_i), .B(
        addresult_12), .C(addresult_13), .Y(\un3_addresult[13] ));
    OA1B \addresult_RNIQKCC[7]  (.A(N_256), .B(\addresult[7]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[7]));
    MX2C un3_addresult_ADD_20x20_slow_I4_un1_CO1_1 (.A(
        ADD_20x20_slow_I1_CO1_m5_i), .B(\addresult_RNIUESN[4]_net_1 ), 
        .S(ADD_20x20_slow_I4_un1_CO1_m11_i), .Y(I4_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        un1_ten_choice_one_0_7_3), .B(\addresult[3]_net_1 ), .C(
        I2_un1_CO1), .Y(\un3_addresult[3] ));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[18]_net_1 ));
    AO18 \addresult_RNIOL9N[4]  (.A(un1_n_s_change_0_1[4]), .B(
        \addresult[4]_net_1 ), .C(d_N_4), .Y(d_N_13));
    OR3B \addresult_RNING0D[19]  (.A(G_1_0_a2_0), .B(
        \addresult[19]_net_1 ), .C(s_addchoice[0]), .Y(N_212));
    XOR3 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        un1_ten_choice_one_0_7_6), .B(\addresult[6]_net_1 ), .C(N236), 
        .Y(\un3_addresult[6] ));
    OA1B \addresult_RNISSCC[9]  (.A(N_256), .B(\addresult[9]_net_1 ), 
        .C(N_33), .Y(signal_data_0_iv_i_0[9]));
    AOI1 \addresult_RNIQBRS7[3]  (.A(signal_data_iv_0_13_3), .B(
        \signal_data_iv_0_12[3] ), .C(signal_data_en[9]), .Y(
        un1_signal_acq_0[3]));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_13));
    AX1E un3_addresult_ADD_20x20_slow_I1_S_0_0 (.A(
        \addresult[0]_net_1 ), .B(un1_ten_choice_one_0_7_0), .C(
        \addresult[1]_net_1 ), .Y(ADD_20x20_slow_I1_S_0_0));
    MIN3 \addresult_RNIIUB24[11]  (.A(I10_un1_CO1), .B(
        \addresult[11]_net_1 ), .C(un1_ten_choice_one_0_7_11), .Y(
        r_N_7_2_i));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[9]_net_1 ));
    DFN1E1C0 \addresult[19]  (.D(\addresult_RNO[19]_net_1 ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .E(
        ADD_20x20_slow_I19_Y_0_m6_e), .Q(\addresult[19]_net_1 ));
    AO18 un3_addresult_ADD_20x20_slow_I1_CO1_m5_i_0 (.A(
        ADD_20x20_slow_I1_CO1tt_m1_e), .B(un1_n_s_change_0_1[1]), .C(
        \addresult[1]_net_1 ), .Y(ADD_20x20_slow_I1_CO1_m5_i_0));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[0]_net_1 ));
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0_7_7), .B(\addresult[7]_net_1 ), .C(
        I6_un1_CO1), .Y(\un3_addresult[7] ));
    NOR3C \addresult_RNI8HEG3[2]  (.A(signal_data_iv_0_1_2), .B(
        \signal_data_iv_0_0[2] ), .C(signal_data_iv_0_9_2), .Y(
        \signal_data_iv_0_12[2] ));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_7_9), .B(\addresult[9]_net_1 ), .C(
        I8_un1_CO1), .Y(\un3_addresult[9] ));
    XOR3 un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        ADD_20x20_slow_I1_CO1_m5_i), .B(\addresult[2]_net_1 ), .C(
        un1_ten_choice_one_0_7_2), .Y(\un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult[1]_net_1 ));
    
endmodule


module add_reg_add_reg_2(
       addresult_RNI5DQA,
       addresult_RNI7DQA,
       addresult_5_10,
       addresult_5_8,
       addresult_RNIDU3E,
       signal_data_0_iv_i_3,
       signal_data_iv_0_0_10,
       signal_data_iv_0_10_0,
       signal_data_iv_0_10_3,
       signal_data_iv_0_10_2,
       un1_ten_choice_one_0_2_0,
       un1_ten_choice_one_0_2_2,
       un1_ten_choice_one_0_2_3,
       un1_ten_choice_one_0_2_4,
       un1_ten_choice_one_0_2_5,
       un1_ten_choice_one_0_2_7,
       un1_ten_choice_one_0_2_8,
       un1_ten_choice_one_0_2_9,
       un1_ten_choice_one_0_2_10,
       un1_ten_choice_one_0_2_6,
       un1_n_s_change_0_1,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_249,
       N_252,
       N_249_0,
       N_215,
       N_210,
       N_192,
       N_189,
       N_179,
       N_147,
       N_139,
       N_131,
       N_123,
       N_155,
       N_171,
       N_251,
       N_241,
       N_238,
       N_208,
       N_205,
       N_224_0,
       N_259,
       N_221,
       N_224
    );
output [12:12] addresult_RNI5DQA;
output [14:14] addresult_RNI7DQA;
output addresult_5_10;
output addresult_5_8;
input  [4:4] addresult_RNIDU3E;
output [11:4] signal_data_0_iv_i_3;
output [1:1] signal_data_iv_0_0_10;
output signal_data_iv_0_10_0;
output signal_data_iv_0_10_3;
output signal_data_iv_0_10_2;
input  un1_ten_choice_one_0_2_0;
input  un1_ten_choice_one_0_2_2;
input  un1_ten_choice_one_0_2_3;
input  un1_ten_choice_one_0_2_4;
input  un1_ten_choice_one_0_2_5;
input  un1_ten_choice_one_0_2_7;
input  un1_ten_choice_one_0_2_8;
input  un1_ten_choice_one_0_2_9;
input  un1_ten_choice_one_0_2_10;
input  un1_ten_choice_one_0_2_6;
input  [2:0] un1_n_s_change_0_1;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
input  N_249;
input  N_252;
input  N_249_0;
input  N_215;
input  N_210;
input  N_192;
input  N_189;
input  N_179;
input  N_147;
input  N_139;
input  N_131;
input  N_123;
input  N_155;
input  N_171;
input  N_251;
input  N_241;
input  N_238;
input  N_208;
input  N_205;
input  N_224_0;
input  N_259;
input  N_221;
input  N_224;

    wire ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0, 
        ADD_20x20_slow_I2_un1_CO1_N_15, 
        ADD_20x20_slow_I2_un1_CO1_m11_i_o4, \addresult_6[2] , 
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_1, ADD_20x20_slow_I7_S_0_0, 
        \addresult_5[7] , ADD_20x20_slow_I6_un1_CO1_0_tz_0, 
        \addresult_5[5] , I4_un1_CO1, \addresult_6[6] , 
        ADD_20x20_slow_I2_S_0_0, ADD_20x20_slow_I2_un1_CO1_m11_i_0, 
        ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0, 
        ADD_20x20_slow_I2_un1_CO1_N_12, N_222, \signal_data_iv_0_5[2] , 
        N_206, \signal_data_iv_0_5[3] , \addresult_6[3] , N_239, 
        \signal_data_iv_0_0_5[1] , \addresult_6[1] , \addresult_6[11] , 
        \addresult_6[8] , \addresult_5[9] , \addresult_6[10] , 
        \addresult_6[4] , N_190, \signal_data_iv_0_5[0] , 
        \addresult_6[0] , ADD_20x20_slow_I11_S_0, I10_un1_CO1, 
        ADD_20x20_slow_I10_S_0, N244, ADD_20x20_slow_I9_S_0, 
        I8_un1_CO1, ADD_20x20_slow_I8_S_0, N240, ADD_20x20_slow_I7_S_0, 
        I6_un1_CO1, ADD_20x20_slow_I6_S_0, N236, ADD_20x20_slow_I5_S_0, 
        ADD_20x20_slow_I4_S_0, N232, ADD_20x20_slow_I3_S_0, 
        ADD_20x20_slow_I2_un1_CO1_m11_i, ADD_20x20_slow_I1_S_0, 
        I0_un1_CO1, ADD_20x20_slow_I2_S_0, ADD_20x20_slow_I1_CO1_0, 
        I1_un3_CO1, ADD_20x20_slow_I6_un1_CO1_0, 
        ADD_20x20_slow_I5_CO1_0, I6_un5_CO1, N248, N254, 
        \addresult_6[12] , I14_un1_CO1, \addresult_6[14] , 
        ADD_20x20_slow_I12_S_0, ADD_20x20_slow_I13_S_0, 
        ADD_20x20_slow_I14_S_0, ADD_20x20_slow_I15_S_0, 
        \addresult_6[17] , \addresult_6[16] , ADD_20x20_slow_I19_Y_0, 
        N270, \addresult_6[18] , \addresult_6[19] , 
        ADD_20x20_slow_I18_S_0, ADD_20x20_slow_I17_S_0, I16_un1_CO1, 
        ADD_20x20_slow_I16_S_0, ADD_20x20_slow_I0_S_0, GND, VCC, GND_0, 
        VCC_0;
    
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        un1_ten_choice_one_0_2_10), .B(\addresult_6[11] ), .C(
        I10_un1_CO1), .Y(ADD_20x20_slow_I11_S_0));
    DFN1C0 \addresult[12]  (.D(ADD_20x20_slow_I12_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[12] ));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_2_7), .B(\addresult_6[8] ), .C(N240), .Y(
        ADD_20x20_slow_I8_S_0));
    OA1 \addresult_RNIJ7HO[4]  (.A(N_251), .B(\addresult_6[4] ), .C(
        addresult_RNIDU3E[4]), .Y(signal_data_0_iv_i_3[4]));
    DFN1C0 \addresult[10]  (.D(ADD_20x20_slow_I10_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[10] ));
    DFN1C0 \addresult[6]  (.D(ADD_20x20_slow_I6_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[6] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(
        ADD_20x20_slow_I2_un1_CO1_m11_i), .B(\addresult_6[3] ), .C(
        un1_ten_choice_one_0_2_2), .Y(N232));
    DFN1C0 \addresult[8]  (.D(ADD_20x20_slow_I8_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[8] ));
    OA1 \addresult_RNILFHO[5]  (.A(N_251), .B(\addresult_5[5] ), .C(
        N_171), .Y(signal_data_0_iv_i_3[5]));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(
        un1_ten_choice_one_0_2_0), .B(\addresult_6[1] ), .C(I0_un1_CO1)
        , .Y(ADD_20x20_slow_I1_S_0));
    OR3A \addresult_RNIUMAF[17]  (.A(\addresult_6[17] ), .B(N_249_0), 
        .C(N_252), .Y(N_239));
    AOI1B \addresult_RNIC9T11[2]  (.A(\addresult_6[2] ), .B(N_259), .C(
        N_224_0), .Y(\signal_data_iv_0_5[2] ));
    OR2 un3_addresult_ADD_20x20_slow_I1_un3_CO1 (.A(
        un1_n_s_change_0_1[1]), .B(I0_un1_CO1), .Y(I1_un3_CO1));
    AOI1B \addresult_RNIA5T11[1]  (.A(\addresult_6[1] ), .B(N_259), .C(
        N_241), .Y(\signal_data_iv_0_0_5[1] ));
    DFN1C0 \addresult[15]  (.D(ADD_20x20_slow_I15_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_5_10));
    OR2 \addresult_RNI5DQA[12]  (.A(\addresult_6[12] ), .B(N_251), .Y(
        addresult_RNI5DQA[12]));
    VCC VCC_i (.Y(VCC));
    OA1 un3_addresult_ADD_20x20_slow_I5_CO1_0 (.A(I4_un1_CO1), .B(
        \addresult_5[5] ), .C(un1_ten_choice_one_0_2_4), .Y(
        ADD_20x20_slow_I5_CO1_0));
    OR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1tt_m1_e (.A(
        \addresult_6[0] ), .B(un1_n_s_change_0_1[0]), .Y(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_1));
    MIN3 un3_addresult_ADD_20x20_slow_I11_CO1 (.A(I10_un1_CO1), .B(
        \addresult_6[11] ), .C(un1_ten_choice_one_0_2_10), .Y(N248));
    AO1 un3_addresult_ADD_20x20_slow_I5_CO1 (.A(\addresult_5[5] ), .B(
        I4_un1_CO1), .C(ADD_20x20_slow_I5_CO1_0), .Y(N236));
    AO1D un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_0 (.A(
        ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0), .B(
        ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0), .C(
        ADD_20x20_slow_I2_un1_CO1_N_12), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_0));
    OAI1 un3_addresult_ADD_20x20_slow_I6_un1_CO1_0 (.A(
        ADD_20x20_slow_I5_CO1_0), .B(ADD_20x20_slow_I6_un1_CO1_0_tz_0), 
        .C(un1_ten_choice_one_0_2_5), .Y(ADD_20x20_slow_I6_un1_CO1_0));
    OR2 \addresult_RNI7DQA[14]  (.A(\addresult_6[14] ), .B(N_251), .Y(
        addresult_RNI7DQA[14]));
    DFN1C0 \addresult[4]  (.D(ADD_20x20_slow_I4_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[4] ));
    AX1 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(un1_n_s_change_0_1[0]), 
        .B(N_224), .C(\addresult_6[0] ), .Y(ADD_20x20_slow_I0_S_0));
    OR3B un3_addresult_ADD_20x20_slow_I13_CO1 (.A(\addresult_6[12] ), 
        .B(addresult_5_8), .C(N248), .Y(N254));
    DFN1C0 \addresult[16]  (.D(ADD_20x20_slow_I16_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[16] ));
    XOR3 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        un1_ten_choice_one_0_2_4), .B(\addresult_5[5] ), .C(I4_un1_CO1)
        , .Y(ADD_20x20_slow_I5_S_0));
    NOR3C \addresult_RNIODE42[1]  (.A(N_239), .B(N_238), .C(
        \signal_data_iv_0_0_5[1] ), .Y(signal_data_iv_0_0_10[1]));
    AOI1B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0 (.A(
        un1_n_s_change_0_1[1]), .B(ADD_20x20_slow_I2_un1_CO1tt_m1_e_1), 
        .C(\addresult_6[1] ), .Y(ADD_20x20_slow_I2_un1_CO1_m11_i_o3_0));
    XNOR2 un3_addresult_ADD_20x20_slow_I14_S_0 (.A(\addresult_6[14] ), 
        .B(N254), .Y(ADD_20x20_slow_I14_S_0));
    OR2B un3_addresult_ADD_20x20_slow_I6_un5_CO1 (.A(\addresult_6[6] ), 
        .B(N236), .Y(I6_un5_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0_2_3), .B(\addresult_6[4] ), .C(N232), .Y(
        ADD_20x20_slow_I4_S_0));
    XOR2 un3_addresult_ADD_20x20_slow_I18_S_0 (.A(\addresult_6[18] ), 
        .B(N270), .Y(ADD_20x20_slow_I18_S_0));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0 (.A(
        un1_n_s_change_0_1[2]), .B(\addresult_6[2] ), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_12));
    DFN1C0 \addresult[5]  (.D(ADD_20x20_slow_I5_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[5] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_6[8] ), .C(un1_ten_choice_one_0_2_7), .Y(I8_un1_CO1)
        );
    NOR2 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_a3_1 (.A(
        ADD_20x20_slow_I2_un1_CO1tt_m1_e_1), .B(un1_n_s_change_0_1[1]), 
        .Y(ADD_20x20_slow_I2_un1_CO1_N_15));
    AX1C un3_addresult_ADD_20x20_slow_I19_Y_0 (.A(N270), .B(
        \addresult_6[18] ), .C(\addresult_6[19] ), .Y(
        ADD_20x20_slow_I19_Y_0));
    OA1 \addresult_RNINNHO[6]  (.A(N_251), .B(\addresult_6[6] ), .C(
        N_179), .Y(signal_data_0_iv_i_3[6]));
    OA1 \addresult_RNIT1AP[11]  (.A(N_251), .B(\addresult_6[11] ), .C(
        N_155), .Y(signal_data_0_iv_i_3[11]));
    DFN1C0 \addresult[2]  (.D(ADD_20x20_slow_I2_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[2] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult_5[7] ), .C(un1_ten_choice_one_0_2_6), .Y(N240));
    NOR2A un3_addresult_ADD_20x20_slow_I14_un1_CO1 (.A(
        \addresult_6[14] ), .B(N254), .Y(I14_un1_CO1));
    AX1C un3_addresult_ADD_20x20_slow_I16_S_0 (.A(I14_un1_CO1), .B(
        addresult_5_10), .C(\addresult_6[16] ), .Y(
        ADD_20x20_slow_I16_S_0));
    DFN1C0 \addresult[3]  (.D(ADD_20x20_slow_I3_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[3] ));
    XOR2 un3_addresult_ADD_20x20_slow_I17_S_0 (.A(\addresult_6[17] ), 
        .B(I16_un1_CO1), .Y(ADD_20x20_slow_I17_S_0));
    DFN1C0 \addresult[14]  (.D(ADD_20x20_slow_I14_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[14] ));
    AO1B un3_addresult_ADD_20x20_slow_I1_CO1_0 (.A(
        un1_ten_choice_one_0_2_0), .B(I0_un1_CO1), .C(\addresult_6[1] )
        , .Y(ADD_20x20_slow_I1_CO1_0));
    XNOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(\addresult_6[12] ), 
        .B(N248), .Y(ADD_20x20_slow_I12_S_0));
    GND GND_i (.Y(GND));
    NOR3C \addresult_RNISLE42[2]  (.A(N_222), .B(N_221), .C(
        \signal_data_iv_0_5[2] ), .Y(signal_data_iv_0_10_2));
    MAJ3 un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(N232), .B(
        \addresult_6[4] ), .C(un1_ten_choice_one_0_2_3), .Y(I4_un1_CO1)
        );
    NOR3C un3_addresult_ADD_20x20_slow_I16_un1_CO1 (.A(I14_un1_CO1), 
        .B(addresult_5_10), .C(\addresult_6[16] ), .Y(I16_un1_CO1));
    XOR2 un3_addresult_ADD_20x20_slow_I7_S_0_0 (.A(\addresult_5[7] ), 
        .B(un1_ten_choice_one_0_2_6), .Y(ADD_20x20_slow_I7_S_0_0));
    NOR2B un3_addresult_ADD_20x20_slow_I17_CO1 (.A(\addresult_6[17] ), 
        .B(I16_un1_CO1), .Y(N270));
    XOR2 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(addresult_5_10), .B(
        I14_un1_CO1), .Y(ADD_20x20_slow_I15_S_0));
    OA1 \addresult_RNIR1AP[10]  (.A(N_251), .B(\addresult_6[10] ), .C(
        N_147), .Y(signal_data_0_iv_i_3[10]));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult_6[10] ), .C(un1_ten_choice_one_0_2_9), .Y(
        I10_un1_CO1));
    OR3A \addresult_RNIVMAF[18]  (.A(\addresult_6[18] ), .B(N_249), .C(
        N_252), .Y(N_222));
    NOR3 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i (.A(N_210), .B(
        ADD_20x20_slow_I2_un1_CO1_m11_i_0), .C(N_215), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i));
    NOR3C \addresult_RNI0UE42[3]  (.A(N_206), .B(N_205), .C(
        \signal_data_iv_0_5[3] ), .Y(signal_data_iv_0_10_3));
    DFN1C0 \addresult[11]  (.D(ADD_20x20_slow_I11_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[11] ));
    OA1 \addresult_RNIR7IO[8]  (.A(N_251), .B(\addresult_6[8] ), .C(
        N_131), .Y(signal_data_0_iv_i_3[8]));
    DFN1C0 \addresult[17]  (.D(ADD_20x20_slow_I17_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[17] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1), .B(
        \addresult_5[9] ), .C(un1_ten_choice_one_0_2_8), .Y(N244));
    AO1 un3_addresult_ADD_20x20_slow_I6_un1_CO1_0_tz_0 (.A(
        \addresult_5[5] ), .B(I4_un1_CO1), .C(\addresult_6[6] ), .Y(
        ADD_20x20_slow_I6_un1_CO1_0_tz_0));
    AOI1B \addresult_RNI81T11[0]  (.A(\addresult_6[0] ), .B(N_259), .C(
        N_192), .Y(\signal_data_iv_0_5[0] ));
    AX1A un3_addresult_ADD_20x20_slow_I2_S_0_0 (.A(
        un1_n_s_change_0_1[2]), .B(N_224), .C(\addresult_6[2] ), .Y(
        ADD_20x20_slow_I2_S_0_0));
    OA1 \addresult_RNITFIO[9]  (.A(N_251), .B(\addresult_5[9] ), .C(
        N_139), .Y(signal_data_0_iv_i_3[9]));
    OR2B un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(I6_un5_CO1), .B(
        ADD_20x20_slow_I6_un1_CO1_0), .Y(I6_un1_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_2_9), .B(\addresult_6[10] ), .C(N244), .Y(
        ADD_20x20_slow_I10_S_0));
    AOI1B \addresult_RNIEDT11[3]  (.A(\addresult_6[3] ), .B(N_259), .C(
        N_208), .Y(\signal_data_iv_0_5[3] ));
    DFN1C0 \addresult[7]  (.D(ADD_20x20_slow_I7_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[7] ));
    OR3A \addresult_RNITMAF[16]  (.A(\addresult_6[16] ), .B(N_249_0), 
        .C(N_252), .Y(N_190));
    AX1 un3_addresult_ADD_20x20_slow_I13_S_0 (.A(N248), .B(
        \addresult_6[12] ), .C(addresult_5_8), .Y(
        ADD_20x20_slow_I13_S_0));
    XOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        un1_ten_choice_one_0_2_2), .B(\addresult_6[3] ), .C(
        ADD_20x20_slow_I2_un1_CO1_m11_i), .Y(ADD_20x20_slow_I3_S_0));
    DFN1C0 \addresult[18]  (.D(ADD_20x20_slow_I18_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[18] ));
    NOR3C \addresult_RNIK5E42[0]  (.A(N_190), .B(N_189), .C(
        \signal_data_iv_0_5[0] ), .Y(signal_data_iv_0_10_0));
    XOR3 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        un1_ten_choice_one_0_2_5), .B(\addresult_6[6] ), .C(N236), .Y(
        ADD_20x20_slow_I6_S_0));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_o4 (.A(
        \addresult_6[2] ), .B(un1_n_s_change_0_1[2]), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_o4));
    OR2 un3_addresult_ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0_0 (.A(
        ADD_20x20_slow_I2_un1_CO1_N_15), .B(
        ADD_20x20_slow_I2_un1_CO1_m11_i_o4), .Y(
        ADD_20x20_slow_I2_un1_CO1_m11_i_a4_0));
    OA1 \addresult_RNIPVHO[7]  (.A(N_251), .B(\addresult_5[7] ), .C(
        N_123), .Y(signal_data_0_iv_i_3[7]));
    OR3A \addresult_RNI0NAF[19]  (.A(\addresult_6[19] ), .B(N_249), .C(
        N_252), .Y(N_206));
    DFN1C0 \addresult[13]  (.D(ADD_20x20_slow_I13_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        addresult_5_8));
    DFN1C0 \addresult[9]  (.D(ADD_20x20_slow_I9_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_5[9] ));
    DFN1C0 \addresult[19]  (.D(ADD_20x20_slow_I19_Y_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[19] ));
    DFN1C0 \addresult[0]  (.D(ADD_20x20_slow_I0_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[0] ));
    OR3B un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(N_224), .B(
        \addresult_6[0] ), .C(un1_n_s_change_0_1[0]), .Y(I0_un1_CO1));
    XOR2 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        ADD_20x20_slow_I7_S_0_0), .B(I6_un1_CO1), .Y(
        ADD_20x20_slow_I7_S_0));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_2_8), .B(\addresult_5[9] ), .C(I8_un1_CO1)
        , .Y(ADD_20x20_slow_I9_S_0));
    AX1C un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        ADD_20x20_slow_I1_CO1_0), .B(I1_un3_CO1), .C(
        ADD_20x20_slow_I2_S_0_0), .Y(ADD_20x20_slow_I2_S_0));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(ADD_20x20_slow_I1_S_0), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_6[1] ));
    
endmodule


module add_reg_add_reg_2_2(
       addresult_RNIVJME,
       un1_n_s_change_0_1,
       un1_ten_choice_one_0_3_0,
       un1_ten_choice_one_0_3_1,
       un1_ten_choice_one_0_3_3,
       un1_ten_choice_one_0_3_10,
       un1_ten_choice_one_0_3_4,
       un1_ten_choice_one_0_3_6,
       un1_ten_choice_one_0_3_7,
       un1_ten_choice_one_0_3_8,
       un1_ten_choice_one_0_3_9,
       un1_ten_choice_one_0_3_11,
       un1_ten_choice_one_0_3_5,
       s_acq_change_0_s_rst,
       signalclkctrl_0_clk_add,
       N_249,
       N_220,
       N_221,
       N_205,
       N_89,
       N_105,
       N_204,
       N_189,
       N_266,
       N_238,
       N_237,
       N_253,
       N_249_0,
       N_188,
       N_177,
       N_169,
       N_153,
       N_145,
       N_137,
       N_129,
       N_121,
       N_113,
       N_252,
       N_97,
       N_219
    );
output [4:4] addresult_RNIVJME;
input  [2:0] un1_n_s_change_0_1;
input  un1_ten_choice_one_0_3_0;
input  un1_ten_choice_one_0_3_1;
input  un1_ten_choice_one_0_3_3;
input  un1_ten_choice_one_0_3_10;
input  un1_ten_choice_one_0_3_4;
input  un1_ten_choice_one_0_3_6;
input  un1_ten_choice_one_0_3_7;
input  un1_ten_choice_one_0_3_8;
input  un1_ten_choice_one_0_3_9;
input  un1_ten_choice_one_0_3_11;
input  un1_ten_choice_one_0_3_5;
input  s_acq_change_0_s_rst;
input  signalclkctrl_0_clk_add;
input  N_249;
output N_220;
output N_221;
output N_205;
output N_89;
output N_105;
output N_204;
output N_189;
input  N_266;
output N_238;
output N_237;
input  N_253;
input  N_249_0;
output N_188;
output N_177;
output N_169;
output N_153;
output N_145;
output N_137;
output N_129;
output N_121;
output N_113;
input  N_252;
output N_97;
input  N_219;

    wire ADD_20x20_slow_I16_un1_CO1_0, \addresult_3[16] , 
        \addresult_2[15] , ADD_20x20_slow_I14_un1_CO1_0, 
        \addresult_3[14] , ADD_20x20_slow_I13_CO1_s, 
        ADD_20x20_slow_I5_S_0_0, \addresult_3[5] , 
        ADD_20x20_slow_I2_S_0_0, \addresult_3[2] , 
        ADD_20x20_slow_I4_un1_CO1_0_tz_0, \addresult_3[3] , 
        ADD_20x20_slow_I2_un1_CO1_m10_i, \addresult_3[4] , 
        ADD_20x20_slow_I2_un1_CO1_m10_i_a4_0, 
        ADD_20x20_slow_I2_un1_CO1_N_16, ADD_20x20_slow_I19_Y_0_m6_e_3, 
        \addresult_2[13] , \addresult_3[18] , 
        ADD_20x20_slow_I19_Y_0_m6_e_2, \addresult_3[17] , 
        \addresult_3[12] , ADD_20x20_slow_I19_Y_0_m6_e_1, 
        \un3_addresult[11] , \addresult_3[11] , I10_un1_CO1, 
        \un3_addresult[9] , \addresult_3[9] , I8_un1_CO1, 
        \un3_addresult[8] , \addresult_3[8] , N240, \un3_addresult[7] , 
        \addresult_2[7] , I6_un1_CO1, \un3_addresult[6] , 
        \addresult_3[6] , N236, \un3_addresult[5] , I4_un1_CO1, 
        \un3_addresult[4] , N232, \un3_addresult[10] , 
        \addresult_3[10] , N244, \un3_addresult[3] , 
        \un3_addresult[2] , ADD_20x20_slow_I1_CO1_0, I1_un3_CO1, 
        \un3_addresult[1] , \addresult_3[1] , I0_un1_CO1, 
        ADD_20x20_slow_I2_un1_CO1_N_11, 
        ADD_20x20_slow_I2_un1_CO1_m10_i_o3_0_tz, 
        ADD_20x20_slow_I2_un1_CO1_N_12, ADD_20x20_slow_I19_Y_0_m6_e_0, 
        I14_un1_CO1, r_N_7_1, I16_un1_CO1, \addresult_3[0] , 
        \addresult_RNO_0[19] , \addresult_3[19] , 
        ADD_20x20_slow_I4_un1_CO1_0, ADD_20x20_slow_I3_CO1_0, 
        I4_un5_CO1, \un3_addresult[12] , \un3_addresult[13] , 
        \un3_addresult[14] , \un3_addresult[15] , \un3_addresult[18] , 
        \un3_addresult[17] , \un3_addresult[0] , \un3_addresult[16] , 
        GND, VCC, GND_0, VCC_0;
    
    NOR2B un3_addresult_ADD_20x20_slow_I13_CO1_s (.A(\addresult_2[13] )
        , .B(\addresult_3[12] ), .Y(ADD_20x20_slow_I13_CO1_s));
    XOR3 un3_addresult_ADD_20x20_slow_I11_S_0 (.A(
        un1_ten_choice_one_0_3_11), .B(\addresult_3[11] ), .C(
        I10_un1_CO1), .Y(\un3_addresult[11] ));
    DFN1C0 \addresult[12]  (.D(\un3_addresult[12] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[12] ));
    XOR3 un3_addresult_ADD_20x20_slow_I8_S_0 (.A(
        un1_ten_choice_one_0_3_8), .B(\addresult_3[8] ), .C(N240), .Y(
        \un3_addresult[8] ));
    OR3A \addresult_RNIAFLB[18]  (.A(\addresult_3[18] ), .B(N_249), .C(
        N_253), .Y(N_220));
    OR2 \addresult_RNI1SME[6]  (.A(\addresult_3[6] ), .B(N_252), .Y(
        N_177));
    OR2 \addresult_RNI34NE[8]  (.A(\addresult_3[8] ), .B(N_252), .Y(
        N_129));
    DFN1C0 \addresult[10]  (.D(\un3_addresult[10] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[10] ));
    DFN1C0 \addresult[6]  (.D(\un3_addresult[6] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[6] ));
    AO1 un3_addresult_ADD_20x20_slow_I3_CO1 (.A(\addresult_3[3] ), .B(
        ADD_20x20_slow_I2_un1_CO1_m10_i), .C(ADD_20x20_slow_I3_CO1_0), 
        .Y(N232));
    MAJ3 \addresult_RNILOOCE[11]  (.A(I10_un1_CO1), .B(
        \addresult_3[11] ), .C(un1_ten_choice_one_0_3_11), .Y(r_N_7_1));
    DFN1C0 \addresult[8]  (.D(\un3_addresult[8] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[8] ));
    XOR3 un3_addresult_ADD_20x20_slow_I1_S_0 (.A(
        un1_ten_choice_one_0_3_1), .B(\addresult_3[1] ), .C(I0_un1_CO1)
        , .Y(\un3_addresult[1] ));
    OR2A un3_addresult_ADD_20x20_slow_I1_un3_CO1 (.A(I0_un1_CO1), .B(
        un1_n_s_change_0_1[1]), .Y(I1_un3_CO1));
    DFN1C0 \addresult[15]  (.D(\un3_addresult[15] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[15] ));
    OA1B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i_a4 (.A(
        ADD_20x20_slow_I2_un1_CO1_m10_i_o3_0_tz), .B(
        un1_n_s_change_0_1[1]), .C(
        ADD_20x20_slow_I2_un1_CO1_m10_i_a4_0), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_11));
    XOR2 \addresult_RNO[19]  (.A(r_N_7_1), .B(\addresult_3[19] ), .Y(
        \addresult_RNO_0[19] ));
    OR3A \addresult_RNIBFLB[19]  (.A(\addresult_3[19] ), .B(N_249_0), 
        .C(N_253), .Y(N_204));
    OR2 \addresult_RNI0OME[5]  (.A(\addresult_3[5] ), .B(N_252), .Y(
        N_169));
    NOR3A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i (.A(N_219), .B(
        ADD_20x20_slow_I2_un1_CO1_N_11), .C(
        ADD_20x20_slow_I2_un1_CO1_N_12), .Y(
        ADD_20x20_slow_I2_un1_CO1_m10_i));
    VCC VCC_i (.Y(VCC));
    MAJ3 un3_addresult_ADD_20x20_slow_I5_CO1 (.A(I4_un1_CO1), .B(
        \addresult_3[5] ), .C(un1_ten_choice_one_0_3_5), .Y(N236));
    OR2 \addresult_RNIVJME[4]  (.A(\addresult_3[4] ), .B(N_252), .Y(
        addresult_RNIVJME[4]));
    DFN1C0 \addresult[4]  (.D(\un3_addresult[4] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[4] ));
    XOR2 un3_addresult_ADD_20x20_slow_I0_S_0 (.A(
        un1_ten_choice_one_0_3_0), .B(\addresult_3[0] ), .Y(
        \un3_addresult[0] ));
    OR2 \addresult_RNIE557[10]  (.A(\addresult_3[10] ), .B(N_252), .Y(
        N_145));
    DFN1C0 \addresult[16]  (.D(\un3_addresult[16] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[16] ));
    XOR2 un3_addresult_ADD_20x20_slow_I5_S_0 (.A(
        ADD_20x20_slow_I5_S_0_0), .B(I4_un1_CO1), .Y(
        \un3_addresult[5] ));
    OR2 \addresult_RNI48NE[9]  (.A(\addresult_3[9] ), .B(N_252), .Y(
        N_137));
    OR3A \addresult_RNI9FLB[17]  (.A(\addresult_3[17] ), .B(N_249_0), 
        .C(N_253), .Y(N_237));
    AX1C un3_addresult_ADD_20x20_slow_I14_S_0 (.A(
        ADD_20x20_slow_I13_CO1_s), .B(r_N_7_1), .C(\addresult_3[14] ), 
        .Y(\un3_addresult[14] ));
    XOR3 un3_addresult_ADD_20x20_slow_I4_S_0 (.A(
        un1_ten_choice_one_0_3_4), .B(\addresult_3[4] ), .C(N232), .Y(
        \un3_addresult[4] ));
    AX1C un3_addresult_ADD_20x20_slow_I18_S_0 (.A(I16_un1_CO1), .B(
        \addresult_3[17] ), .C(\addresult_3[18] ), .Y(
        \un3_addresult[18] ));
    DFN1C0 \addresult[5]  (.D(\un3_addresult[5] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[5] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I8_un1_CO1 (.A(N240), .B(
        \addresult_3[8] ), .C(un1_ten_choice_one_0_3_8), .Y(I8_un1_CO1)
        );
    DFN1C0 \addresult[2]  (.D(\un3_addresult[2] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[2] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        \addresult_2[7] ), .C(un1_ten_choice_one_0_3_7), .Y(N240));
    NOR2B un3_addresult_ADD_20x20_slow_I14_un1_CO1 (.A(
        ADD_20x20_slow_I14_un1_CO1_0), .B(r_N_7_1), .Y(I14_un1_CO1));
    AO1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0_tz_0 (.A(
        \addresult_3[3] ), .B(ADD_20x20_slow_I2_un1_CO1_m10_i), .C(
        \addresult_3[4] ), .Y(ADD_20x20_slow_I4_un1_CO1_0_tz_0));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e (.A(
        ADD_20x20_slow_I19_Y_0_m6_e_2), .B(
        ADD_20x20_slow_I19_Y_0_m6_e_1), .C(
        ADD_20x20_slow_I19_Y_0_m6_e_3), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_0));
    OR2B \addresult_RNIIP6J[3]  (.A(\addresult_3[3] ), .B(N_266), .Y(
        N_205));
    AX1C un3_addresult_ADD_20x20_slow_I16_S_0 (.A(I14_un1_CO1), .B(
        \addresult_2[15] ), .C(\addresult_3[16] ), .Y(
        \un3_addresult[16] ));
    DFN1C0 \addresult[3]  (.D(\un3_addresult[3] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[3] ));
    XOR2 un3_addresult_ADD_20x20_slow_I17_S_0 (.A(\addresult_3[17] ), 
        .B(I16_un1_CO1), .Y(\un3_addresult[17] ));
    AO1A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i_a4_0_0 (.A(
        un1_n_s_change_0_1[2]), .B(\addresult_3[2] ), .C(
        ADD_20x20_slow_I2_un1_CO1_N_16), .Y(
        ADD_20x20_slow_I2_un1_CO1_m10_i_a4_0));
    DFN1C0 \addresult[14]  (.D(\un3_addresult[14] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[14] ));
    OAI1 un3_addresult_ADD_20x20_slow_I1_CO1_0 (.A(I0_un1_CO1), .B(
        un1_ten_choice_one_0_3_1), .C(\addresult_3[1] ), .Y(
        ADD_20x20_slow_I1_CO1_0));
    XOR2 un3_addresult_ADD_20x20_slow_I12_S_0 (.A(r_N_7_1), .B(
        \addresult_3[12] ), .Y(\un3_addresult[12] ));
    GND GND_i (.Y(GND));
    OR2 un3_addresult_ADD_20x20_slow_I4_un1_CO1 (.A(I4_un5_CO1), .B(
        ADD_20x20_slow_I4_un1_CO1_0), .Y(I4_un1_CO1));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_1 (.A(
        \addresult_3[14] ), .B(\addresult_3[16] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_1));
    NOR2B un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_2 (.A(
        \addresult_3[17] ), .B(\addresult_3[12] ), .Y(
        ADD_20x20_slow_I19_Y_0_m6_e_2));
    NOR2B un3_addresult_ADD_20x20_slow_I16_un1_CO1 (.A(
        ADD_20x20_slow_I16_un1_CO1_0), .B(I14_un1_CO1), .Y(I16_un1_CO1)
        );
    OR2 \addresult_RNIH557[13]  (.A(\addresult_2[13] ), .B(N_252), .Y(
        N_97));
    XOR2 un3_addresult_ADD_20x20_slow_I15_S_0 (.A(\addresult_2[15] ), 
        .B(I14_un1_CO1), .Y(\un3_addresult[15] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I10_un1_CO1 (.A(N244), .B(
        \addresult_3[10] ), .C(un1_ten_choice_one_0_3_10), .Y(
        I10_un1_CO1));
    DFN1C0 \addresult[11]  (.D(\un3_addresult[11] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[11] ));
    OR3A \addresult_RNI8FLB[16]  (.A(\addresult_3[16] ), .B(N_249_0), 
        .C(N_253), .Y(N_188));
    OA1 un3_addresult_ADD_20x20_slow_I4_un1_CO1_0 (.A(
        ADD_20x20_slow_I3_CO1_0), .B(ADD_20x20_slow_I4_un1_CO1_0_tz_0), 
        .C(un1_ten_choice_one_0_3_4), .Y(ADD_20x20_slow_I4_un1_CO1_0));
    OR2 \addresult_RNI20NE[7]  (.A(\addresult_2[7] ), .B(N_252), .Y(
        N_121));
    DFN1C0 \addresult[17]  (.D(\un3_addresult[17] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[17] ));
    MAJ3 un3_addresult_ADD_20x20_slow_I9_CO1 (.A(I8_un1_CO1), .B(
        \addresult_3[9] ), .C(un1_ten_choice_one_0_3_9), .Y(N244));
    AX1A un3_addresult_ADD_20x20_slow_I2_S_0_0 (.A(
        un1_n_s_change_0_1[2]), .B(N_219), .C(\addresult_3[2] ), .Y(
        ADD_20x20_slow_I2_S_0_0));
    OA1C un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i_o3_0_tz (.A(
        \addresult_3[0] ), .B(un1_n_s_change_0_1[0]), .C(
        \addresult_3[1] ), .Y(ADD_20x20_slow_I2_un1_CO1_m10_i_o3_0_tz));
    MAJ3 un3_addresult_ADD_20x20_slow_I6_un1_CO1 (.A(N236), .B(
        \addresult_3[6] ), .C(un1_ten_choice_one_0_3_6), .Y(I6_un1_CO1)
        );
    XOR2 un3_addresult_ADD_20x20_slow_I5_S_0_0 (.A(\addresult_3[5] ), 
        .B(un1_ten_choice_one_0_3_5), .Y(ADD_20x20_slow_I5_S_0_0));
    NOR2B un3_addresult_ADD_20x20_slow_I4_un5_CO1 (.A(\addresult_3[4] )
        , .B(N232), .Y(I4_un5_CO1));
    XOR3 un3_addresult_ADD_20x20_slow_I10_S_0 (.A(
        un1_ten_choice_one_0_3_10), .B(\addresult_3[10] ), .C(N244), 
        .Y(\un3_addresult[10] ));
    OR2 \addresult_RNIJ557[15]  (.A(\addresult_2[15] ), .B(N_252), .Y(
        N_113));
    DFN1C0 \addresult[7]  (.D(\un3_addresult[7] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[7] ));
    NOR3C un3_addresult_ADD_20x20_slow_I19_Y_0_m6_e_3 (.A(
        \addresult_2[13] ), .B(\addresult_3[18] ), .C(
        \addresult_2[15] ), .Y(ADD_20x20_slow_I19_Y_0_m6_e_3));
    OR2B \addresult_RNIFD6J[0]  (.A(\addresult_3[0] ), .B(N_266), .Y(
        N_189));
    AX1C un3_addresult_ADD_20x20_slow_I13_S_0 (.A(\addresult_3[12] ), 
        .B(r_N_7_1), .C(\addresult_2[13] ), .Y(\un3_addresult[13] ));
    XOR3 un3_addresult_ADD_20x20_slow_I3_S_0 (.A(
        un1_ten_choice_one_0_3_3), .B(\addresult_3[3] ), .C(
        ADD_20x20_slow_I2_un1_CO1_m10_i), .Y(\un3_addresult[3] ));
    OR2 \addresult_RNIG557[12]  (.A(\addresult_3[12] ), .B(N_252), .Y(
        N_89));
    OR2B \addresult_RNIHL6J[2]  (.A(\addresult_3[2] ), .B(N_266), .Y(
        N_221));
    DFN1C0 \addresult[18]  (.D(\un3_addresult[18] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[18] ));
    NOR2B un3_addresult_ADD_20x20_slow_I16_un1_CO1_0 (.A(
        \addresult_3[16] ), .B(\addresult_2[15] ), .Y(
        ADD_20x20_slow_I16_un1_CO1_0));
    OR2B \addresult_RNIGH6J[1]  (.A(\addresult_3[1] ), .B(N_266), .Y(
        N_238));
    NOR2A un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i_a4_0 (.A(
        un1_n_s_change_0_1[2]), .B(\addresult_3[2] ), .Y(
        ADD_20x20_slow_I2_un1_CO1_N_12));
    XOR3 un3_addresult_ADD_20x20_slow_I6_S_0 (.A(
        un1_ten_choice_one_0_3_6), .B(\addresult_3[6] ), .C(N236), .Y(
        \un3_addresult[6] ));
    NOR3B un3_addresult_ADD_20x20_slow_I2_un1_CO1_m10_i_a3_1 (.A(
        \addresult_3[0] ), .B(\addresult_3[1] ), .C(
        un1_n_s_change_0_1[0]), .Y(ADD_20x20_slow_I2_un1_CO1_N_16));
    DFN1C0 \addresult[13]  (.D(\un3_addresult[13] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_2[13] ));
    NOR2B un3_addresult_ADD_20x20_slow_I14_un1_CO1_0 (.A(
        \addresult_3[14] ), .B(ADD_20x20_slow_I13_CO1_s), .Y(
        ADD_20x20_slow_I14_un1_CO1_0));
    OR2 \addresult_RNII557[14]  (.A(\addresult_3[14] ), .B(N_252), .Y(
        N_105));
    DFN1C0 \addresult[9]  (.D(\un3_addresult[9] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[9] ));
    DFN1E1C0 \addresult[19]  (.D(\addresult_RNO_0[19] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .E(
        ADD_20x20_slow_I19_Y_0_m6_e_0), .Q(\addresult_3[19] ));
    OA1 un3_addresult_ADD_20x20_slow_I3_CO1_0 (.A(
        ADD_20x20_slow_I2_un1_CO1_m10_i), .B(\addresult_3[3] ), .C(
        un1_ten_choice_one_0_3_3), .Y(ADD_20x20_slow_I3_CO1_0));
    OR2 \addresult_RNIF557[11]  (.A(\addresult_3[11] ), .B(N_252), .Y(
        N_153));
    DFN1C0 \addresult[0]  (.D(\un3_addresult[0] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[0] ));
    NOR2B un3_addresult_ADD_20x20_slow_I0_un1_CO1 (.A(
        un1_ten_choice_one_0_3_0), .B(\addresult_3[0] ), .Y(I0_un1_CO1)
        );
    XOR3 un3_addresult_ADD_20x20_slow_I7_S_0 (.A(
        un1_ten_choice_one_0_3_7), .B(\addresult_2[7] ), .C(I6_un1_CO1)
        , .Y(\un3_addresult[7] ));
    XOR3 un3_addresult_ADD_20x20_slow_I9_S_0 (.A(
        un1_ten_choice_one_0_3_9), .B(\addresult_3[9] ), .C(I8_un1_CO1)
        , .Y(\un3_addresult[9] ));
    AX1C un3_addresult_ADD_20x20_slow_I2_S_0 (.A(
        ADD_20x20_slow_I1_CO1_0), .B(I1_un3_CO1), .C(
        ADD_20x20_slow_I2_S_0_0), .Y(\un3_addresult[2] ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1C0 \addresult[1]  (.D(\un3_addresult[1] ), .CLK(
        signalclkctrl_0_clk_add), .CLR(s_acq_change_0_s_rst), .Q(
        \addresult_3[1] ));
    
endmodule


module signalclkctrl(
       s_acqnum,
       s_periodnum,
       s_stripnum,
       s_acq_change_0_s_load_0,
       s_acq_change_0_s_load,
       GLA,
       s_acq_change_0_s_rst,
       signalclkctrl_0_entop,
       signal_acq_0_Signal_acq_clk,
       clkout,
       signalclkctrl_0_clk_add
    );
input  [15:0] s_acqnum;
input  [3:0] s_periodnum;
input  [11:0] s_stripnum;
input  s_acq_change_0_s_load_0;
input  s_acq_change_0_s_load;
input  GLA;
input  s_acq_change_0_s_rst;
output signalclkctrl_0_entop;
output signal_acq_0_Signal_acq_clk;
input  clkout;
output signalclkctrl_0_clk_add;

    wire clk_add_i, N_50, N_42, \DWACT_FINC_E[0] , N_19, 
        \DWACT_FINC_E[4] , N_4, \DWACT_FINC_E[7] , \DWACT_FINC_E[6] , 
        un1_count_NE_11, un1_count_NE_2, un1_count_NE_1, 
        un1_count_NE_7, un1_count_NE_10, \count_RNIHUU33[12]_net_1 , 
        un1_count_11_i, un1_count_NE_5, un1_count_NE_9, un1_count_9_i, 
        un1_count_5_i, un1_count_NE_4, un1_count_0_i, enclk6_NE_8, 
        \count[13]_net_1 , \count[10]_net_1 , un1_count_10_0_0_net_1, 
        un1_count_8_i, \count[7]_net_1 , un1_count_7_0_0_net_1, 
        un1_count_6_i, \count[4]_net_1 , un1_count_4_0_0_net_1, 
        un1_count_3_i, \count[2]_net_1 , un1_count_2_0_0_1, 
        un1_count_1_0_i, enclk6_NE_11, enclk6_NE_2, enclk6_NE_1, 
        enclk6_NE_7, enclk6_NE_10, enclk6_10_i, enclk6_8_i, 
        enclk6_NE_6, enclk6_NE_9, enclk6_NE_3, enclk6_NE_4, enclk6_0_i, 
        \count[11]_net_1 , I_66_0, enclk6_12_i, \count[6]_net_1 , 
        I_31_0, enclk6_7_i, \count[9]_net_1 , I_52_0, enclk6_5_i, 
        \count[3]_net_1 , I_13_1, enclk6_4_i, \count[1]_net_1 , I_5_1, 
        enclk6_2_i, un1_count_3_0_0, \perioddata[3]_net_1 , 
        \perioddata[2]_net_1 , N142, un1_count_1_1_0_0, 
        \perioddata[1]_net_1 , I8_un1_CO1, N152, N146, 
        \perioddata[0]_net_1 , \count[0]_net_1 , I0_un1_CO1, 
        I2_un1_CO1, I4_un1_CO1, \count[5]_net_1 , N160, 
        \count[8]_net_1 , I10_un1_CO1, un1_count_i, enclk6_NE, enclk8, 
        I_115_0, ADD_16x16_slow_I11_S_0, I10_un1_CO1_0, 
        \data[11]_net_1 , ADD_16x16_slow_I10_S_0, N212, 
        \data[10]_net_1 , ADD_16x16_slow_I9_S_0, I8_un1_CO1_0, 
        \data[9]_net_1 , ADD_16x16_slow_I8_S_0, N208, \data[8]_net_1 , 
        ADD_16x16_slow_I7_S_0, I6_un1_CO1, \data[7]_net_1 , 
        ADD_16x16_slow_I6_S_0, N204, \data[6]_net_1 , 
        ADD_16x16_slow_I5_S_0, I4_un1_CO1_0, \data[5]_net_1 , 
        ADD_16x16_slow_I4_S_0, N200, \data[4]_net_1 , 
        ADD_16x16_slow_I3_S_0, I2_un1_CO1_0, \data[3]_net_1 , 
        ADD_16x16_slow_I2_S_0, N196, \data[2]_net_1 , 
        ADD_16x16_slow_I1_S_0, I0_un1_CO1_0, \data[1]_net_1 , N216, 
        \data[0]_net_1 , N222, \data[12]_net_1 , \data[13]_net_1 , 
        ADD_16x16_slow_I0_S_0, ADD_16x16_slow_I12_S_0, 
        ADD_16x16_slow_I13_S_0, ADD_16x16_slow_I14_S_0, 
        \data[14]_net_1 , ADD_16x16_slow_I15_Y_0, \data[15]_net_1 , 
        I_9_1, I_20_1, I_24_1, I_38_1, I_45_0, I_56_0, 
        \count[12]_net_1 , count_c13, count_c12, count_n14, 
        \count[14]_net_1 , count_n15, \count[15]_net_1 , enadd_net_1, 
        enclk_net_1, count_c2, count_c4, count_c6, count_c8, count_c10, 
        entop_RNO_net_1, enadd_RNO_net_1, enclk_RNO_net_1, count_n1, 
        count_n2, count_n3, count_n4, count_n5, count_n6, count_n7, 
        count_n8, count_n9, count_n10, count_n11, count_n12, count_n13, 
        \count_RNO_0[0] , N_9, \DWACT_FINC_E[2] , \DWACT_FINC_E[5] , 
        N_16, \DWACT_FINC_E[3] , N_24, N_29, N_34, \DWACT_FINC_E[1] , 
        N_39, N_47, \DWACT_COMP0_E[1] , \DWACT_COMP0_E[2] , 
        \DWACT_COMP0_E[0] , \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , N_21, N_20, N_19_0, N_16_0, 
        N_18, N_17, N_15, N_12, N_13, N_14, \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \DWACT_BL_EQUAL_0_E[3] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[0] , 
        \DWACT_BL_EQUAL_0_E[1] , \DWACT_BL_EQUAL_0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] , \ACT_LT4_E_0[3] , 
        \ACT_LT4_E_0[6] , \ACT_LT4_E_0[10] , \ACT_LT4_E_0[7] , 
        \ACT_LT4_E_0[8] , \ACT_LT4_E_0[5] , \ACT_LT4_E_0[4] , 
        \ACT_LT4_E_0[0] , \ACT_LT4_E_0[1] , \ACT_LT4_E_0[2] , 
        \ACT_LT3_E[3] , \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , 
        \ACT_LT3_E[1] , \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E_0[2] , 
        \DWACT_BL_EQUAL_0_E_0[1] , \DWACT_BL_EQUAL_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E[6] , \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] , 
        \DWACT_BL_EQUAL_0_E_0[3] , \DWACT_BL_EQUAL_0_E[4] , 
        \DWACT_BL_EQUAL_0_E[5] , \DWACT_BL_EQUAL_0_E_1[0] , 
        \DWACT_BL_EQUAL_0_E_1[1] , \DWACT_BL_EQUAL_0_E_1[2] , GND, VCC, 
        GND_0, VCC_0;
    
    OR2B enclk_RNI44A5 (.A(enclk_net_1), .B(clkout), .Y(
        signal_acq_0_Signal_acq_clk));
    MAJ3 un1_data_ADD_16x16_slow_I10_un1_CO1 (.A(N212), .B(
        s_stripnum[10]), .C(\data[10]_net_1 ), .Y(I10_un1_CO1_0));
    XA1 \count_RNII7U44[4]  (.A(\count[4]_net_1 ), .B(
        un1_count_4_0_0_net_1), .C(un1_count_3_i), .Y(un1_count_NE_2));
    XOR2 un1_stripnum_I_20 (.A(N_42), .B(s_stripnum[4]), .Y(I_20_1));
    DFN1E1 \data[5]  (.D(s_acqnum[5]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[5]_net_1 ));
    DFN1E1C0 \count[15]  (.D(count_n15), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[15]_net_1 ));
    NOR2A un1_count_1_0_I_76 (.A(ADD_16x16_slow_I5_S_0), .B(
        \count[5]_net_1 ), .Y(\ACT_LT4_E[0] ));
    AX1 \count_RNO[6]  (.A(count_c4), .B(\count[5]_net_1 ), .C(
        \count[6]_net_1 ), .Y(count_n6));
    DFN1C0 enclk (.D(enclk_RNO_net_1), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .Q(enclk_net_1));
    AND3 un1_stripnum_I_62 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[5] ), .Y(
        \DWACT_FINC_E[6] ));
    XA1A \count_RNI5E2H4[11]  (.A(\count[11]_net_1 ), .B(I_66_0), .C(
        enclk6_12_i), .Y(enclk6_NE_6));
    XNOR2 \count_RNO[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_n3));
    XOR2 un1_stripnum_I_5 (.A(s_stripnum[0]), .B(s_stripnum[1]), .Y(
        I_5_1));
    AX1E un1_count_10_0_0 (.A(I8_un1_CO1), .B(s_stripnum[9]), .C(
        s_stripnum[10]), .Y(un1_count_10_0_0_net_1));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[9]_net_1 ));
    XOR2 un1_data_ADD_16x16_slow_I14_S_0 (.A(N222), .B(
        \data[14]_net_1 ), .Y(ADD_16x16_slow_I14_S_0));
    NOR2A un1_count_1_0_I_47 (.A(\count[11]_net_1 ), .B(
        ADD_16x16_slow_I11_S_0), .Y(\ACT_LT4_E_0[7] ));
    AO1C un1_count_1_0_I_101 (.A(\count[3]_net_1 ), .B(
        ADD_16x16_slow_I3_S_0), .C(N_15), .Y(N_20));
    OR3B \count_RNIQVK71[4]  (.A(\count[3]_net_1 ), .B(
        \count[4]_net_1 ), .C(count_c2), .Y(count_c4));
    XA1A \count_RNIG0MK2[2]  (.A(\count[2]_net_1 ), .B(
        un1_count_2_0_0_1), .C(un1_count_1_0_i), .Y(un1_count_NE_1));
    XOR3 \count_RNI9JL13[8]  (.A(N160), .B(s_stripnum[8]), .C(
        \count[8]_net_1 ), .Y(un1_count_8_i));
    DFN1E1 \data[9]  (.D(s_acqnum[9]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[9]_net_1 ));
    XNOR2 \count_RNIBO9V1[7]  (.A(I_38_1), .B(\count[7]_net_1 ), .Y(
        enclk6_7_i));
    DFN1E1 \data[10]  (.D(s_acqnum[10]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[10]_net_1 ));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[8]_net_1 ));
    OA1A un1_count_1_0_I_102 (.A(N_16_0), .B(N_18), .C(N_17), .Y(N_21));
    XOR2 \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .Y(count_n1));
    XOR3 un1_data_ADD_16x16_slow_I8_S_0 (.A(N208), .B(\data[8]_net_1 ), 
        .C(s_stripnum[8]), .Y(ADD_16x16_slow_I8_S_0));
    AX1 \count_RNO[12]  (.A(count_c10), .B(\count[11]_net_1 ), .C(
        \count[12]_net_1 ), .Y(count_n12));
    XNOR2 \count_RNI16GA1[4]  (.A(I_20_1), .B(\count[4]_net_1 ), .Y(
        enclk6_4_i));
    NOR3C un1_stripnum_1_0_0_ADD_12x12_slow_I10_un1_CO1 (.A(I8_un1_CO1)
        , .B(s_stripnum[9]), .C(s_stripnum[10]), .Y(I10_un1_CO1));
    MAJ3 un1_data_ADD_16x16_slow_I5_CO1 (.A(I4_un1_CO1_0), .B(
        s_stripnum[5]), .C(\data[5]_net_1 ), .Y(N204));
    XNOR2 un1_count_1_0_I_5 (.A(\count[13]_net_1 ), .B(
        ADD_16x16_slow_I13_S_0), .Y(\DWACT_BL_EQUAL_0_E[4] ));
    DFN1E1 \data[13]  (.D(s_acqnum[13]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[13]_net_1 ));
    XOR2 \perioddata_RNI7POD[3]  (.A(\perioddata[3]_net_1 ), .B(
        s_stripnum[3]), .Y(un1_count_3_0_0));
    DFN1C0 enadd (.D(enadd_RNO_net_1), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .Q(enadd_net_1));
    XOR3 un1_data_ADD_16x16_slow_I6_S_0 (.A(N204), .B(\data[6]_net_1 ), 
        .C(s_stripnum[6]), .Y(ADD_16x16_slow_I6_S_0));
    AO1C un1_count_1_0_I_99 (.A(\count[2]_net_1 ), .B(
        ADD_16x16_slow_I2_S_0), .C(N_12), .Y(N_18));
    AX1C \count_RNO[2]  (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(count_n2));
    NOR2A un1_count_1_0_I_81 (.A(ADD_16x16_slow_I8_S_0), .B(
        \count[8]_net_1 ), .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_count_1_0_I_65 (.A(\count[8]_net_1 ), .B(
        ADD_16x16_slow_I8_S_0), .Y(\DWACT_BL_EQUAL_0_E[3] ));
    XNOR2 \count_RNO[11]  (.A(count_c10), .B(\count[11]_net_1 ), .Y(
        count_n11));
    XNOR2 \count_RNIA3LS[2]  (.A(I_9_1), .B(\count[2]_net_1 ), .Y(
        enclk6_2_i));
    OR2A un1_count_1_0_I_48 (.A(\count[12]_net_1 ), .B(
        ADD_16x16_slow_I12_S_0), .Y(\ACT_LT4_E_0[8] ));
    NOR2B un1_stripnum_I_72 (.A(\DWACT_FINC_E[7] ), .B(
        \DWACT_FINC_E[6] ), .Y(N_4));
    XNOR2 un1_count_1_0_I_21 (.A(\count[15]_net_1 ), .B(
        ADD_16x16_slow_I15_Y_0), .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    XOR2 un1_stripnum_I_31 (.A(N_34), .B(s_stripnum[6]), .Y(I_31_0));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[10]_net_1 ));
    XNOR2 \count_RNIQJA72[10]  (.A(I_56_0), .B(\count[10]_net_1 ), .Y(
        enclk6_10_i));
    OR2A un1_count_1_0_I_31 (.A(ADD_16x16_slow_I15_Y_0), .B(
        \count[15]_net_1 ), .Y(\ACT_LT3_E[4] ));
    AO1 un1_count_1_0_I_110 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), 
        .B(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(\DWACT_COMP0_E[2] ));
    DFN1E1 \data[4]  (.D(s_acqnum[4]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[4]_net_1 ));
    XNOR3 \count_RNI3A0V1[3]  (.A(I2_un1_CO1), .B(un1_count_3_0_0), .C(
        \count[3]_net_1 ), .Y(un1_count_3_i));
    XOR2 un1_stripnum_I_9 (.A(N_50), .B(s_stripnum[2]), .Y(I_9_1));
    DFN1E1 \data[11]  (.D(s_acqnum[11]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[11]_net_1 ));
    NOR2A un1_stripnum_1_0_0_ADD_12x12_slow_I4_un1_CO1 (.A(
        s_stripnum[4]), .B(N146), .Y(I4_un1_CO1));
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[5]_net_1 ));
    AND3 un1_stripnum_I_34 (.A(s_stripnum[3]), .B(s_stripnum[4]), .C(
        s_stripnum[5]), .Y(\DWACT_FINC_E[2] ));
    NOR3C \count_RNIQTKU8[10]  (.A(enclk6_10_i), .B(enclk6_8_i), .C(
        enclk6_NE_6), .Y(enclk6_NE_10));
    OR2 un1_stripnum_1_0_0_ADD_12x12_slow_I0_un1_CO1 (.A(s_stripnum[0])
        , .B(\perioddata[0]_net_1 ), .Y(I0_un1_CO1));
    XA1A \count_RNI30HE5[7]  (.A(\count[7]_net_1 ), .B(
        un1_count_7_0_0_net_1), .C(un1_count_6_i), .Y(un1_count_NE_4));
    OR3B \count_RNIL10PH5[10]  (.A(enclk6_NE), .B(un1_count_i), .C(
        I_115_0), .Y(enclk8));
    NOR3C \count_RNIIRBCC[10]  (.A(\count_RNIHUU33[12]_net_1 ), .B(
        un1_count_11_i), .C(un1_count_NE_5), .Y(un1_count_NE_10));
    XNOR2 un1_count_1_0_I_6 (.A(\count[14]_net_1 ), .B(
        ADD_16x16_slow_I14_S_0), .Y(\DWACT_BL_EQUAL_0_E[5] ));
    NOR3C un1_data_ADD_16x16_slow_I13_CO1 (.A(\data[12]_net_1 ), .B(
        N216), .C(\data[13]_net_1 ), .Y(N222));
    XNOR2 un1_count_1_0_I_63 (.A(\count[6]_net_1 ), .B(
        ADD_16x16_slow_I6_S_0), .Y(\DWACT_BL_EQUAL_0_E[1] ));
    AND2A un1_count_1_0_I_29 (.A(ADD_16x16_slow_I14_S_0), .B(
        \count[14]_net_1 ), .Y(\ACT_LT3_E[2] ));
    NOR3B \count_RNI0OBO[13]  (.A(un1_count_0_i), .B(enclk6_NE_8), .C(
        \count[13]_net_1 ), .Y(un1_count_NE_7));
    AND3 un1_stripnum_I_37 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(s_stripnum[6]), .Y(N_29));
    AND3 un1_count_1_0_I_66 (.A(\DWACT_BL_EQUAL_0_E[0] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    NOR2A \count_RNINGVI2[13]  (.A(\count[13]_net_1 ), .B(count_c12), 
        .Y(count_c13));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[4]_net_1 ));
    AND3 un1_stripnum_I_55 (.A(\DWACT_FINC_E[4] ), .B(s_stripnum[8]), 
        .C(s_stripnum[9]), .Y(N_16));
    GND GND_i (.Y(GND));
    NOR3B \count_RNI6AGH[13]  (.A(enclk6_0_i), .B(enclk6_NE_8), .C(
        \count[13]_net_1 ), .Y(enclk6_NE_7));
    DFN1E1C0 \count[12]  (.D(count_n12), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[12]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1P0 \count[0]  (.D(\count_RNO_0[0] ), .CLK(clkout), .PRE(
        s_acq_change_0_s_rst), .Q(\count[0]_net_1 ));
    NOR2A un1_count_1_0_I_95 (.A(ADD_16x16_slow_I0_S_0), .B(
        \count[0]_net_1 ), .Y(N_14));
    XOR3 un1_data_ADD_16x16_slow_I9_S_0 (.A(I8_un1_CO1_0), .B(
        \data[9]_net_1 ), .C(s_stripnum[9]), .Y(ADD_16x16_slow_I9_S_0));
    AX1C un1_data_ADD_16x16_slow_I13_S_0 (.A(\data[12]_net_1 ), .B(
        N216), .C(\data[13]_net_1 ), .Y(ADD_16x16_slow_I13_S_0));
    XNOR2 \count_RNIRR762[8]  (.A(I_45_0), .B(\count[8]_net_1 ), .Y(
        enclk6_8_i));
    DFN1E1 \perioddata[2]  (.D(s_periodnum[2]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\perioddata[2]_net_1 ));
    XOR3 \count_RNIAGPJ2[6]  (.A(N152), .B(s_stripnum[6]), .C(
        \count[6]_net_1 ), .Y(un1_count_6_i));
    XNOR2 \count_RNO[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_n5));
    MAJ3 un1_data_ADD_16x16_slow_I9_CO1 (.A(I8_un1_CO1_0), .B(
        s_stripnum[9]), .C(\data[9]_net_1 ), .Y(N212));
    DFN1E1 \data[1]  (.D(s_acqnum[1]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[1]_net_1 ));
    MAJ3 un1_data_ADD_16x16_slow_I3_CO1 (.A(I2_un1_CO1_0), .B(
        s_stripnum[3]), .C(\data[3]_net_1 ), .Y(N200));
    AX1C \count_RNO[15]  (.A(\count[14]_net_1 ), .B(count_c13), .C(
        \count[15]_net_1 ), .Y(count_n15));
    AND3 un1_stripnum_I_69 (.A(s_stripnum[9]), .B(s_stripnum[10]), .C(
        s_stripnum[11]), .Y(\DWACT_FINC_E[7] ));
    AOI1A un1_count_1_0_I_50 (.A(\ACT_LT4_E_0[3] ), .B(
        \ACT_LT4_E_0[6] ), .C(\ACT_LT4_E_0[10] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ));
    DFN1E1 \data[6]  (.D(s_acqnum[6]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[6]_net_1 ));
    OR3B \count_RNI5FHN1[5]  (.A(\count[5]_net_1 ), .B(
        \count[6]_net_1 ), .C(count_c4), .Y(count_c6));
    AND3 un1_stripnum_I_12 (.A(s_stripnum[0]), .B(s_stripnum[1]), .C(
        s_stripnum[2]), .Y(N_47));
    XOR2 un1_stripnum_I_13 (.A(N_47), .B(s_stripnum[3]), .Y(I_13_1));
    AND3 un1_count_1_0_I_9 (.A(\DWACT_BL_EQUAL_0_E_0[3] ), .B(
        \DWACT_BL_EQUAL_0_E[4] ), .C(\DWACT_BL_EQUAL_0_E[5] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    AOI1A un1_count_1_0_I_85 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), 
        .C(\ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    OR2A un1_count_1_0_I_77 (.A(ADD_16x16_slow_I6_S_0), .B(
        \count[6]_net_1 ), .Y(\ACT_LT4_E[1] ));
    OR2A un1_count_1_0_I_93 (.A(ADD_16x16_slow_I1_S_0), .B(
        \count[1]_net_1 ), .Y(N_12));
    DFN1E1 \perioddata[3]  (.D(s_periodnum[3]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\perioddata[3]_net_1 ));
    XOR2 un1_data_ADD_16x16_slow_I12_S_0 (.A(N216), .B(
        \data[12]_net_1 ), .Y(ADD_16x16_slow_I12_S_0));
    DFN1E1 \data[8]  (.D(s_acqnum[8]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[8]_net_1 ));
    DFN1E1 \perioddata[1]  (.D(s_periodnum[1]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\perioddata[1]_net_1 ));
    XNOR3 \count_RNISKRC2[5]  (.A(I4_un1_CO1), .B(s_stripnum[5]), .C(
        \count[5]_net_1 ), .Y(un1_count_5_i));
    NOR2B un1_data_ADD_16x16_slow_I0_un1_CO1 (.A(s_stripnum[0]), .B(
        \data[0]_net_1 ), .Y(I0_un1_CO1_0));
    XOR3 un1_data_ADD_16x16_slow_I2_S_0 (.A(N196), .B(\data[2]_net_1 ), 
        .C(s_stripnum[2]), .Y(ADD_16x16_slow_I2_S_0));
    XOR3 \perioddata_RNI9J991[2]  (.A(s_stripnum[2]), .B(
        \perioddata[2]_net_1 ), .C(N142), .Y(un1_count_2_0_0_1));
    VCC VCC_i (.Y(VCC));
    OR2A un1_count_1_0_I_41 (.A(ADD_16x16_slow_I10_S_0), .B(
        \count[10]_net_1 ), .Y(\ACT_LT4_E_0[1] ));
    XNOR3 \count_RNILJE31[1]  (.A(I0_un1_CO1), .B(un1_count_1_1_0_0), 
        .C(\count[1]_net_1 ), .Y(un1_count_1_0_i));
    AND3 un1_stripnum_I_30 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[1] ), .C(s_stripnum[5]), .Y(N_34));
    XOR3 un1_data_ADD_16x16_slow_I7_S_0 (.A(I6_un1_CO1), .B(
        \data[7]_net_1 ), .C(s_stripnum[7]), .Y(ADD_16x16_slow_I7_S_0));
    OR2A un1_count_1_0_I_96 (.A(ADD_16x16_slow_I4_S_0), .B(
        \count[4]_net_1 ), .Y(N_15));
    XOR2 \count_RNO[14]  (.A(count_c13), .B(\count[14]_net_1 ), .Y(
        count_n14));
    XOR2 un1_count_4_0_0 (.A(s_stripnum[4]), .B(N146), .Y(
        un1_count_4_0_0_net_1));
    XNOR2 un1_count_1_0_I_62 (.A(\count[5]_net_1 ), .B(
        ADD_16x16_slow_I5_S_0), .Y(\DWACT_BL_EQUAL_0_E[0] ));
    AO1 un1_count_1_0_I_115 (.A(\DWACT_COMP0_E[1] ), .B(
        \DWACT_COMP0_E[2] ), .C(\DWACT_COMP0_E[0] ), .Y(I_115_0));
    XA1A \count_RNIQ0KU3[9]  (.A(\count[9]_net_1 ), .B(I_52_0), .C(
        enclk6_5_i), .Y(enclk6_NE_3));
    DFN1E1C0 \count[13]  (.D(count_n13), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[13]_net_1 ));
    MAJ3 un1_data_ADD_16x16_slow_I2_un1_CO1 (.A(N196), .B(
        s_stripnum[2]), .C(\data[2]_net_1 ), .Y(I2_un1_CO1_0));
    AND3 un1_count_1_0_I_8 (.A(\DWACT_BL_EQUAL_0_E_1[0] ), .B(
        \DWACT_BL_EQUAL_0_E_1[1] ), .C(\DWACT_BL_EQUAL_0_E_1[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ));
    NOR2A un1_count_1_0_I_83 (.A(\count[7]_net_1 ), .B(
        ADD_16x16_slow_I7_S_0), .Y(\ACT_LT4_E[7] ));
    XNOR2 un1_count_1_0_I_2 (.A(\count[10]_net_1 ), .B(
        ADD_16x16_slow_I10_S_0), .Y(\DWACT_BL_EQUAL_0_E_1[1] ));
    DFN1E1 \data[7]  (.D(s_acqnum[7]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[7]_net_1 ));
    AOI1A un1_count_1_0_I_49 (.A(\ACT_LT4_E_0[7] ), .B(
        \ACT_LT4_E_0[8] ), .C(\ACT_LT4_E_0[5] ), .Y(\ACT_LT4_E_0[10] ));
    XOR2 un1_stripnum_I_66 (.A(N_9), .B(s_stripnum[11]), .Y(I_66_0));
    XOR2 un1_stripnum_I_52 (.A(N_19), .B(s_stripnum[9]), .Y(I_52_0));
    XNOR2 un1_count_1_0_I_64 (.A(\count[7]_net_1 ), .B(
        ADD_16x16_slow_I7_S_0), .Y(\DWACT_BL_EQUAL_0_E[2] ));
    DFN1E1 \data[14]  (.D(s_acqnum[14]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[14]_net_1 ));
    XNOR2 un1_count_1_0_I_3 (.A(\count[15]_net_1 ), .B(
        ADD_16x16_slow_I15_Y_0), .Y(\DWACT_BL_EQUAL_0_E[6] ));
    AND2A un1_count_1_0_I_78 (.A(ADD_16x16_slow_I6_S_0), .B(
        \count[6]_net_1 ), .Y(\ACT_LT4_E[2] ));
    XOR2 \count_RNO[0]  (.A(enclk8), .B(\count[0]_net_1 ), .Y(
        \count_RNO_0[0] ));
    DFN1E1 \data[0]  (.D(s_acqnum[0]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[0]_net_1 ));
    OR3B \count_RNIJT2I2[12]  (.A(\count[11]_net_1 ), .B(
        \count[12]_net_1 ), .C(count_c10), .Y(count_c12));
    AOI1A un1_count_1_0_I_86 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), 
        .C(\ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    AOI1A un1_count_1_0_I_33 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), 
        .C(\ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ));
    NOR2B un1_stripnum_I_51 (.A(s_stripnum[8]), .B(\DWACT_FINC_E[4] ), 
        .Y(N_19));
    AO1 un1_count_1_0_I_57 (.A(\DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ), .B(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[0] ), .Y(\DWACT_COMP0_E[0] ));
    XA1A \count_RNI7HLN3[6]  (.A(\count[6]_net_1 ), .B(I_31_0), .C(
        enclk6_7_i), .Y(enclk6_NE_4));
    XOR3 un1_data_ADD_16x16_slow_I4_S_0 (.A(N200), .B(\data[4]_net_1 ), 
        .C(s_stripnum[4]), .Y(ADD_16x16_slow_I4_S_0));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[1]_net_1 ));
    XNOR2 \count_RNO[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_n7));
    NOR2 \count_RNIB6P1[15]  (.A(\count[15]_net_1 ), .B(
        \count[14]_net_1 ), .Y(enclk6_NE_8));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[3]_net_1 ));
    XNOR2 \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_n9));
    DFN1E1 \data[15]  (.D(s_acqnum[15]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[15]_net_1 ));
    OR2A enclk_RNO (.A(enclk6_NE), .B(enclk_net_1), .Y(enclk_RNO_net_1)
        );
    MAJ3 un1_data_ADD_16x16_slow_I4_un1_CO1 (.A(N200), .B(
        s_stripnum[4]), .C(\data[4]_net_1 ), .Y(I4_un1_CO1_0));
    XNOR2 un1_count_1_0_I_19 (.A(\count[13]_net_1 ), .B(
        ADD_16x16_slow_I13_S_0), .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    XOR3 \perioddata_RNIHULL[0]  (.A(s_stripnum[0]), .B(
        \perioddata[0]_net_1 ), .C(\count[0]_net_1 ), .Y(un1_count_0_i)
        );
    AND2 un1_count_1_0_I_67 (.A(\DWACT_BL_EQUAL_0_E[3] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    OA1 un1_count_1_0_I_103 (.A(N_21), .B(N_20), .C(N_19_0), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    MAJ3 un1_data_ADD_16x16_slow_I6_un1_CO1 (.A(N204), .B(
        s_stripnum[6]), .C(\data[6]_net_1 ), .Y(I6_un1_CO1));
    OR2B un1_stripnum_1_0_0_ADD_12x12_slow_I5_CO1 (.A(s_stripnum[5]), 
        .B(I4_un1_CO1), .Y(N152));
    NOR3C \count_RNIPF04B[5]  (.A(un1_count_9_i), .B(un1_count_5_i), 
        .C(un1_count_NE_4), .Y(un1_count_NE_9));
    OR2A un1_count_1_0_I_94 (.A(\count[2]_net_1 ), .B(
        ADD_16x16_slow_I2_S_0), .Y(N_13));
    NOR2A un1_count_1_0_I_45 (.A(ADD_16x16_slow_I12_S_0), .B(
        \count[12]_net_1 ), .Y(\ACT_LT4_E_0[5] ));
    AX1 \count_RNO[4]  (.A(count_c2), .B(\count[3]_net_1 ), .C(
        \count[4]_net_1 ), .Y(count_n4));
    NOR2A un1_stripnum_1_0_0_ADD_12x12_slow_I8_un1_CO1 (.A(
        s_stripnum[8]), .B(N160), .Y(I8_un1_CO1));
    XNOR2 \count_RNO[13]  (.A(count_c12), .B(\count[13]_net_1 ), .Y(
        count_n13));
    NOR2B un1_stripnum_I_19 (.A(s_stripnum[3]), .B(\DWACT_FINC_E[0] ), 
        .Y(N_42));
    NOR2A un1_count_1_0_I_82 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), 
        .Y(\ACT_LT4_E[6] ));
    XNOR3 \count_RNIGUU33[11]  (.A(I10_un1_CO1), .B(s_stripnum[11]), 
        .C(\count[11]_net_1 ), .Y(un1_count_11_i));
    OR2A un1_count_1_0_I_80 (.A(ADD_16x16_slow_I7_S_0), .B(
        \count[7]_net_1 ), .Y(\ACT_LT4_E[4] ));
    MAJ3 un1_data_ADD_16x16_slow_I8_un1_CO1 (.A(N208), .B(
        s_stripnum[8]), .C(\data[8]_net_1 ), .Y(I8_un1_CO1_0));
    AND3 un1_count_1_0_I_22 (.A(\DWACT_BL_EQUAL_0_E_0[2] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_0[0] ), .Y(
        \DWACT_CMPLE_PO0_DWACT_COMP0_E[1] ));
    XOR2 \perioddata_RNI3HOD[1]  (.A(\perioddata[1]_net_1 ), .B(
        s_stripnum[1]), .Y(un1_count_1_1_0_0));
    AND2A un1_count_1_0_I_32 (.A(ADD_16x16_slow_I15_Y_0), .B(
        \count[15]_net_1 ), .Y(\ACT_LT3_E[5] ));
    DFN1E1 \data[2]  (.D(s_acqnum[2]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[2]_net_1 ));
    XNOR2 un1_count_1_0_I_20 (.A(\count[14]_net_1 ), .B(
        ADD_16x16_slow_I14_S_0), .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    XNOR2 \count_RNI37H82[12]  (.A(N_4), .B(\count[12]_net_1 ), .Y(
        enclk6_12_i));
    XOR2 un1_stripnum_I_45 (.A(N_24), .B(s_stripnum[8]), .Y(I_45_0));
    AOI1A un1_count_1_0_I_30 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), 
        .C(\ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    AND3 un1_stripnum_I_48 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(
        \DWACT_FINC_E[4] ));
    OR2A un1_count_1_0_I_100 (.A(\count[4]_net_1 ), .B(
        ADD_16x16_slow_I4_S_0), .Y(N_19_0));
    GND GND_i_0 (.Y(GND_0));
    NOR2B enadd_RNIFR95 (.A(enadd_net_1), .B(clkout), .Y(clk_add_i));
    OR2A un1_count_1_0_I_84 (.A(\count[8]_net_1 ), .B(
        ADD_16x16_slow_I8_S_0), .Y(\ACT_LT4_E[8] ));
    XNOR2 un1_count_1_0_I_4 (.A(\count[11]_net_1 ), .B(
        ADD_16x16_slow_I11_S_0), .Y(\DWACT_BL_EQUAL_0_E_1[2] ));
    AOI1A un1_count_1_0_I_43 (.A(\ACT_LT4_E_0[0] ), .B(
        \ACT_LT4_E_0[1] ), .C(\ACT_LT4_E_0[2] ), .Y(\ACT_LT4_E_0[3] ));
    OR3C \count_RNIJ0PN[2]  (.A(\count[0]_net_1 ), .B(\count[1]_net_1 )
        , .C(\count[2]_net_1 ), .Y(count_c2));
    NOR3C \count_RNI200I7[13]  (.A(un1_count_NE_2), .B(un1_count_NE_1), 
        .C(un1_count_NE_7), .Y(un1_count_NE_11));
    MAJ3 un1_data_ADD_16x16_slow_I7_CO1 (.A(I6_un1_CO1), .B(
        s_stripnum[7]), .C(\data[7]_net_1 ), .Y(N208));
    XNOR2 \count_RNIETDH1[5]  (.A(I_24_1), .B(\count[5]_net_1 ), .Y(
        enclk6_5_i));
    AO1A enadd_RNO (.A(un1_count_i), .B(enclk6_NE), .C(enadd_net_1), 
        .Y(enadd_RNO_net_1));
    NOR2A un1_count_1_0_I_46 (.A(\ACT_LT4_E_0[4] ), .B(
        \ACT_LT4_E_0[5] ), .Y(\ACT_LT4_E_0[6] ));
    XOR2 \count_RNINGQE[0]  (.A(s_stripnum[0]), .B(\count[0]_net_1 ), 
        .Y(enclk6_0_i));
    NOR2B entop_RNO (.A(signalclkctrl_0_entop), .B(enclk8), .Y(
        entop_RNO_net_1));
    AO1C un1_count_1_0_I_97 (.A(ADD_16x16_slow_I1_S_0), .B(
        \count[1]_net_1 ), .C(N_14), .Y(N_16_0));
    AND3 un1_stripnum_I_59 (.A(s_stripnum[6]), .B(s_stripnum[7]), .C(
        s_stripnum[8]), .Y(\DWACT_FINC_E[5] ));
    AX1E \count_RNIHUU33[12]  (.A(I10_un1_CO1), .B(s_stripnum[11]), .C(
        \count[12]_net_1 ), .Y(\count_RNIHUU33[12]_net_1 ));
    MAJ3 un1_data_ADD_16x16_slow_I1_CO1 (.A(I0_un1_CO1_0), .B(
        s_stripnum[1]), .C(\data[1]_net_1 ), .Y(N196));
    XNOR3 \count_RNIQQJ83[9]  (.A(I8_un1_CO1), .B(s_stripnum[9]), .C(
        \count[9]_net_1 ), .Y(un1_count_9_i));
    MAJ3 un1_data_ADD_16x16_slow_I11_CO1 (.A(I10_un1_CO1_0), .B(
        s_stripnum[11]), .C(\data[11]_net_1 ), .Y(N216));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[7]_net_1 ));
    AND3 un1_stripnum_I_16 (.A(s_stripnum[0]), .B(s_stripnum[1]), .C(
        s_stripnum[2]), .Y(\DWACT_FINC_E[0] ));
    OR3B \count_RNIKEE72[8]  (.A(\count[7]_net_1 ), .B(
        \count[8]_net_1 ), .C(count_c6), .Y(count_c8));
    AOI1A un1_count_1_0_I_79 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), 
        .C(\ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    XNOR2 un1_count_1_0_I_1 (.A(\count[9]_net_1 ), .B(
        ADD_16x16_slow_I9_S_0), .Y(\DWACT_BL_EQUAL_0_E_1[0] ));
    DFN1P0 entop (.D(entop_RNO_net_1), .CLK(clkout), .PRE(
        s_acq_change_0_s_rst), .Q(signalclkctrl_0_entop));
    AND3 un1_stripnum_I_23 (.A(\DWACT_FINC_E[0] ), .B(s_stripnum[3]), 
        .C(s_stripnum[4]), .Y(N_39));
    MIN3 un1_stripnum_1_0_0_ADD_12x12_slow_I3_CO1 (.A(I2_un1_CO1), .B(
        s_stripnum[3]), .C(\perioddata[3]_net_1 ), .Y(N146));
    MAJ3 un1_stripnum_1_0_0_ADD_12x12_slow_I1_CO1 (.A(I0_un1_CO1), .B(
        s_stripnum[1]), .C(\perioddata[1]_net_1 ), .Y(N142));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[6]_net_1 ));
    XOR3 un1_data_ADD_16x16_slow_I5_S_0 (.A(I4_un1_CO1_0), .B(
        \data[5]_net_1 ), .C(s_stripnum[5]), .Y(ADD_16x16_slow_I5_S_0));
    NOR2A un1_count_1_0_I_27 (.A(ADD_16x16_slow_I13_S_0), .B(
        \count[13]_net_1 ), .Y(\ACT_LT3_E[0] ));
    AX1C un1_data_ADD_16x16_slow_I15_Y_0 (.A(\data[14]_net_1 ), .B(
        N222), .C(\data[15]_net_1 ), .Y(ADD_16x16_slow_I15_Y_0));
    XOR2 un1_stripnum_I_24 (.A(N_39), .B(s_stripnum[5]), .Y(I_24_1));
    OA1A un1_count_1_0_I_98 (.A(\count[3]_net_1 ), .B(
        ADD_16x16_slow_I3_S_0), .C(N_13), .Y(N_17));
    XOR3 un1_data_ADD_16x16_slow_I1_S_0 (.A(I0_un1_CO1_0), .B(
        \data[1]_net_1 ), .C(s_stripnum[1]), .Y(ADD_16x16_slow_I1_S_0));
    XA1A \count_RNIMO2E2[3]  (.A(\count[3]_net_1 ), .B(I_13_1), .C(
        enclk6_4_i), .Y(enclk6_NE_2));
    CLKINT enadd_RNIFR95_0 (.A(clk_add_i), .Y(signalclkctrl_0_clk_add));
    AND3 un1_stripnum_I_65 (.A(\DWACT_FINC_E[6] ), .B(s_stripnum[9]), 
        .C(s_stripnum[10]), .Y(N_9));
    XOR3 un1_data_ADD_16x16_slow_I3_S_0 (.A(I2_un1_CO1_0), .B(
        \data[3]_net_1 ), .C(s_stripnum[3]), .Y(ADD_16x16_slow_I3_S_0));
    MAJ3 un1_stripnum_1_0_0_ADD_12x12_slow_I2_un1_CO1 (.A(N142), .B(
        s_stripnum[2]), .C(\perioddata[2]_net_1 ), .Y(I2_un1_CO1));
    AND2 un1_stripnum_I_27 (.A(s_stripnum[3]), .B(s_stripnum[4]), .Y(
        \DWACT_FINC_E[1] ));
    XOR2 un1_stripnum_I_56 (.A(N_16), .B(s_stripnum[10]), .Y(I_56_0));
    AND2A un1_count_1_0_I_42 (.A(ADD_16x16_slow_I10_S_0), .B(
        \count[10]_net_1 ), .Y(\ACT_LT4_E_0[2] ));
    AX1 un1_count_7_0_0 (.A(N152), .B(s_stripnum[6]), .C(s_stripnum[7])
        , .Y(un1_count_7_0_0_net_1));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[2]_net_1 ));
    NOR2A un1_count_1_0_I_40 (.A(ADD_16x16_slow_I9_S_0), .B(
        \count[9]_net_1 ), .Y(\ACT_LT4_E_0[0] ));
    AND2 un1_stripnum_I_41 (.A(s_stripnum[6]), .B(s_stripnum[7]), .Y(
        \DWACT_FINC_E[3] ));
    NOR3C \count_RNI6UVH4[13]  (.A(enclk6_NE_2), .B(enclk6_NE_1), .C(
        enclk6_NE_7), .Y(enclk6_NE_11));
    AX1 \count_RNO[8]  (.A(count_c6), .B(\count[7]_net_1 ), .C(
        \count[8]_net_1 ), .Y(count_n8));
    OR3C \count_RNI1EU6L[10]  (.A(enclk6_NE_10), .B(enclk6_NE_9), .C(
        enclk6_NE_11), .Y(enclk6_NE));
    DFN1E1 \perioddata[0]  (.D(s_periodnum[0]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\perioddata[0]_net_1 ));
    XOR2 un1_data_ADD_16x16_slow_I0_S_0 (.A(s_stripnum[0]), .B(
        \data[0]_net_1 ), .Y(ADD_16x16_slow_I0_S_0));
    OR3B un1_stripnum_1_0_0_ADD_12x12_slow_I7_CO1 (.A(s_stripnum[6]), 
        .B(s_stripnum[7]), .C(N152), .Y(N160));
    XOR3 un1_data_ADD_16x16_slow_I10_S_0 (.A(N212), .B(
        \data[10]_net_1 ), .C(s_stripnum[10]), .Y(
        ADD_16x16_slow_I10_S_0));
    OR2A un1_count_1_0_I_28 (.A(ADD_16x16_slow_I14_S_0), .B(
        \count[14]_net_1 ), .Y(\ACT_LT3_E[1] ));
    AND3 un1_stripnum_I_44 (.A(\DWACT_FINC_E[0] ), .B(
        \DWACT_FINC_E[2] ), .C(\DWACT_FINC_E[3] ), .Y(N_24));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[11]_net_1 ));
    OR2A un1_count_1_0_I_44 (.A(ADD_16x16_slow_I11_S_0), .B(
        \count[11]_net_1 ), .Y(\ACT_LT4_E_0[4] ));
    XA1A \count_RNIARCI1[1]  (.A(\count[1]_net_1 ), .B(I_5_1), .C(
        enclk6_2_i), .Y(enclk6_NE_1));
    NOR2B \count_RNI1I9M7[6]  (.A(enclk6_NE_3), .B(enclk6_NE_4), .Y(
        enclk6_NE_9));
    XOR2 un1_stripnum_I_38 (.A(N_29), .B(s_stripnum[7]), .Y(I_38_1));
    DFN1E1 \data[12]  (.D(s_acqnum[12]), .CLK(GLA), .E(
        s_acq_change_0_s_load_0), .Q(\data[12]_net_1 ));
    DFN1E1C0 \count[14]  (.D(count_n14), .CLK(clkout), .CLR(
        s_acq_change_0_s_rst), .E(enclk8), .Q(\count[14]_net_1 ));
    AX1 \count_RNO[10]  (.A(count_c8), .B(\count[9]_net_1 ), .C(
        \count[10]_net_1 ), .Y(count_n10));
    XA1 \count_RNIHUD46[10]  (.A(\count[10]_net_1 ), .B(
        un1_count_10_0_0_net_1), .C(un1_count_8_i), .Y(un1_count_NE_5));
    OR3B \count_RNIEN9G2[10]  (.A(\count[9]_net_1 ), .B(
        \count[10]_net_1 ), .C(count_c8), .Y(count_c10));
    AND3 un1_count_1_0_I_10 (.A(\DWACT_BL_EQUAL_0_E[6] ), .B(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), .C(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E_0[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    XOR3 un1_data_ADD_16x16_slow_I11_S_0 (.A(I10_un1_CO1_0), .B(
        \data[11]_net_1 ), .C(s_stripnum[11]), .Y(
        ADD_16x16_slow_I11_S_0));
    OR3C \count_RNIDBC2V[10]  (.A(un1_count_NE_10), .B(un1_count_NE_9), 
        .C(un1_count_NE_11), .Y(un1_count_i));
    XNOR2 un1_count_1_0_I_7 (.A(\count[12]_net_1 ), .B(
        ADD_16x16_slow_I12_S_0), .Y(\DWACT_BL_EQUAL_0_E_0[3] ));
    NOR2B un1_stripnum_I_8 (.A(s_stripnum[1]), .B(s_stripnum[0]), .Y(
        N_50));
    DFN1E1 \data[3]  (.D(s_acqnum[3]), .CLK(GLA), .E(
        s_acq_change_0_s_load), .Q(\data[3]_net_1 ));
    
endmodule


module signal_acq(
       un1_add_reg_4_i_0,
       un1_add_reg_4_i_2,
       ADC_c,
       addresult_0_0,
       addresult_0_2,
       addresult_RNIJE5C,
       addresult,
       un1_signal_acq_0,
       addresult_4_0,
       addresult_4_2,
       addresult_RNI8MQ7,
       s_stripnum,
       s_periodnum,
       s_acqnum,
       un1_n_s_change_0_1,
       addresult_5_0,
       addresult_5_2,
       addresult_RNI7DQA,
       addresult_RNI5DQA,
       s_addchoice,
       top_code_0_n_s_ctrl_0,
       N_104,
       N_88,
       N_86,
       N_27_i_0,
       N_22_i_0,
       N_18_i_0,
       N_16_i_0,
       N_14_i_0,
       N_12_i_0,
       N_20_i_0,
       N_25_i_0,
       N_92,
       N_108,
       N_99,
       N_115,
       N_107,
       N_91,
       N_97,
       N_113,
       N_105,
       N_89,
       N_87,
       N_95,
       N_111,
       signal_acq_0_Signal_acq_clk,
       GLA,
       s_acq_change_0_s_load,
       s_acq_change_0_s_load_0,
       scan_scale_sw_0_s_start,
       ddsclkout_c,
       s_acq_change_0_s_rst,
       N_33,
       N_256,
       N_255,
       N_253,
       N_251,
       N_39
    );
output un1_add_reg_4_i_0;
output un1_add_reg_4_i_2;
input  [2:0] ADC_c;
output addresult_0_0;
output addresult_0_2;
output [14:14] addresult_RNIJE5C;
output [15:12] addresult;
output [3:0] un1_signal_acq_0;
output addresult_4_0;
output addresult_4_2;
output [14:14] addresult_RNI8MQ7;
input  [11:0] s_stripnum;
input  [3:0] s_periodnum;
input  [15:0] s_acqnum;
input  [11:0] un1_n_s_change_0_1;
output addresult_5_0;
output addresult_5_2;
output [14:14] addresult_RNI7DQA;
output [12:12] addresult_RNI5DQA;
input  [4:0] s_addchoice;
input  top_code_0_n_s_ctrl_0;
output N_104;
output N_88;
output N_86;
output N_27_i_0;
output N_22_i_0;
output N_18_i_0;
output N_16_i_0;
output N_14_i_0;
output N_12_i_0;
output N_20_i_0;
output N_25_i_0;
output N_92;
output N_108;
output N_99;
output N_115;
output N_107;
output N_91;
output N_97;
output N_113;
output N_105;
output N_89;
output N_87;
output N_95;
output N_111;
output signal_acq_0_Signal_acq_clk;
input  GLA;
input  s_acq_change_0_s_load;
input  s_acq_change_0_s_load_0;
input  scan_scale_sw_0_s_start;
input  ddsclkout_c;
input  s_acq_change_0_s_rst;
output N_33;
output N_256;
output N_255;
output N_253;
output N_251;
output N_39;

    wire N_249_0, G_1_0_a2_0_net_1, \signal_data_en[9] , N_249, N_250, 
        N_252, N_254, N_262, N_267, N_273, N_271, N_270, N_266, N_263, 
        N_259, \addresult_RNIDU3E[4] , \signal_data_0_iv_i_3[4] , 
        \signal_data_0_iv_i_3[5] , \signal_data_0_iv_i_3[6] , 
        \signal_data_0_iv_i_3[7] , \signal_data_0_iv_i_3[8] , 
        \signal_data_0_iv_i_3[9] , \signal_data_0_iv_i_3[10] , 
        \signal_data_0_iv_i_3[11] , \signal_data_iv_0_0_10[1] , 
        \signal_data_iv_0_10[0] , \signal_data_iv_0_10[3] , 
        \signal_data_iv_0_10[2] , \un1_ten_choice_one_0_2[1] , 
        \un1_ten_choice_one_0_2[3] , \un1_ten_choice_one_0_2[4] , 
        \un1_ten_choice_one_0_2[5] , \un1_ten_choice_one_0_2[6] , 
        \un1_ten_choice_one_0_2[8] , \un1_ten_choice_one_0_2[9] , 
        \un1_ten_choice_one_0_2[10] , \un1_ten_choice_one_0_2[11] , 
        \un1_ten_choice_one_0_2[7] , signalclkctrl_0_clk_add, N_215, 
        N_210, N_192, N_189, N_179, N_147, N_139, N_131, N_123, N_155, 
        N_171, N_241, N_238, N_208, N_205, N_224, N_221, N_224_0, 
        clkout, signalclkctrl_0_entop, \addresult_RNIFE5C[10] , 
        \signal_data_0_iv_i_2[4] , \signal_data_0_iv_i_2[5] , 
        \signal_data_0_iv_i_2[6] , \signal_data_0_iv_i_2[7] , 
        \signal_data_0_iv_i_2[8] , \signal_data_0_iv_i_2[9] , 
        \signal_data_0_iv_i_2[10] , \signal_data_0_iv_i_2[11] , 
        \addresult_RNIBOIB[5] , \signal_data_0_iv_i_5[4] , 
        \signal_data_0_iv_i_5[5] , \signal_data_0_iv_i_5[6] , 
        \signal_data_0_iv_i_5[7] , \signal_data_0_iv_i_5[8] , 
        \signal_data_0_iv_i_5[9] , \signal_data_0_iv_i_5[10] , 
        \signal_data_0_iv_i_5[11] , \signal_data_iv_0_0_3[1] , 
        \signal_data_iv_0_0_9[1] , \signal_data_iv_0_3[0] , 
        \signal_data_iv_0_3[3] , \signal_data_iv_0_3[2] , 
        \signal_data_iv_0_9[0] , \signal_data_iv_0_9[3] , 
        \signal_data_iv_0_9[2] , \un1_ten_choice_one_0_5[0] , 
        \un1_ten_choice_one_0_5[1] , \un1_ten_choice_one_0_5[2] , 
        \un1_ten_choice_one_0_5[3] , \un1_ten_choice_one_0_5[4] , 
        \un1_ten_choice_one_0_5[5] , \un1_ten_choice_one_0_5[6] , 
        \un1_ten_choice_one_0_5[7] , \un1_ten_choice_one_0_5[8] , 
        \un1_ten_choice_one_0_5[9] , \un1_ten_choice_one_0_5[10] , 
        \un1_ten_choice_one_0_5[11] , N_216, N_184, N_200, N_233, 
        N_214, N_186, N_174, N_158, N_134, N_126, N_118, N_150, N_235, 
        N_202, N_218, N_223, \addresult_RNIVJME[4] , 
        \un1_ten_choice_one_0_3[0] , \un1_ten_choice_one_0_3[1] , 
        \un1_ten_choice_one_0_3[3] , \un1_ten_choice_one_0_3[10] , 
        \un1_ten_choice_one_0_3[4] , \un1_ten_choice_one_0_3[6] , 
        \un1_ten_choice_one_0_3[7] , \un1_ten_choice_one_0_3[8] , 
        \un1_ten_choice_one_0_3[9] , \un1_ten_choice_one_0_3[11] , 
        \un1_ten_choice_one_0_3[5] , N_220, N_204, N_237, N_188, N_177, 
        N_169, N_153, N_145, N_137, N_129, N_121, N_219, 
        \signal_data_iv_0_0_6[1] , \signal_data_iv_0_6[0] , 
        \signal_data_iv_0_6[3] , \signal_data_iv_0_6[2] , 
        \un1_ten_choice_one_0_1[0] , \un1_ten_choice_one_0_1[2] , 
        \un1_ten_choice_one_0_1[10] , \un1_ten_choice_one_0_1[5] , 
        \un1_ten_choice_one_0_1[9] , \un1_ten_choice_one_0_1[7] , 
        \un1_ten_choice_one_0_1[1] , \un1_ten_choice_one_0_1[8] , 
        \un1_ten_choice_one_0_1[4] , \un1_ten_choice_one_0_1[6] , 
        \un1_ten_choice_one_0_1[11] , N_194, N_243, N_210_0, N_226, 
        N_213, N_216_0, \signal_data_0_iv_i_0[4] , 
        \signal_data_0_iv_i_0[5] , \signal_data_0_iv_i_0[6] , 
        \signal_data_0_iv_i_0[7] , \signal_data_0_iv_i_0[8] , 
        \signal_data_0_iv_i_0[9] , \signal_data_0_iv_i_0[10] , 
        \signal_data_0_iv_i_0[11] , \signal_data_iv_0_0_13[1] , 
        \signal_data_iv_0_13[0] , \signal_data_iv_0_13[3] , 
        \signal_data_iv_0_13[2] , \un1_ten_choice_one_0[0] , 
        \un1_ten_choice_one_0[1] , \un1_ten_choice_one_0[2] , 
        \un1_ten_choice_one_0[3] , \un1_ten_choice_one_0[4] , 
        \un1_ten_choice_one_0[5] , \un1_ten_choice_one_0[6] , 
        \un1_ten_choice_one_0[7] , \un1_ten_choice_one_0[8] , 
        \un1_ten_choice_one_0[9] , \un1_ten_choice_one_0[10] , 
        \un1_ten_choice_one_0[11] , N_222, N_196, N_245, N_212, N_228, 
        \addrout[0] , \addrout[1] , \addrout[2] , \addrout[3] , 
        \dataeight_0_a2_0_0[0] , \signal_data_iv_0_0_1[1] , 
        \signal_data_iv_0_1[0] , \signal_data_iv_0_1[3] , 
        \signal_data_iv_0_1[2] , \un1_ten_choice_one_0_7[2] , 
        \un1_ten_choice_one_0_7[3] , \un1_ten_choice_one_0_7[5] , 
        \un1_ten_choice_one_0_7[6] , \un1_ten_choice_one_0_7[7] , 
        \un1_ten_choice_one_0_7[8] , \un1_ten_choice_one_0_7[9] , 
        \un1_ten_choice_one_0_7[10] , \un1_ten_choice_one_0_7[11] , 
        \un1_ten_choice_one_0_7[0] , N_182, N_231, N_198, N_214_0, 
        N_220_0, \un1_ten_choice_one_0_6[1] , 
        \un1_ten_choice_one_0_6[2] , \un1_ten_choice_one_0_6[3] , 
        \un1_ten_choice_one_0_6[4] , \un1_ten_choice_one_0_6[5] , 
        \un1_ten_choice_one_0_6[6] , \un1_ten_choice_one_0_6[7] , 
        \un1_ten_choice_one_0_6[8] , \un1_ten_choice_one_0_6[9] , 
        \un1_ten_choice_one_0_6[10] , \un1_ten_choice_one_0_6[11] , 
        N_221_0, N_212_0, \un1_ten_choice_one_0_4[0] , 
        \un1_ten_choice_one_0_4[3] , \un1_ten_choice_one_0_4[1] , 
        \un1_ten_choice_one_0_4[4] , \un1_ten_choice_one_0_4[5] , 
        \un1_ten_choice_one_0_4[7] , \un1_ten_choice_one_0_4[8] , 
        \un1_ten_choice_one_0_4[9] , \un1_ten_choice_one_0_4[10] , 
        \un1_ten_choice_one_0_4[11] , \un1_ten_choice_one_0_4[6] , 
        N_211, N_217, GND, VCC, GND_0, VCC_0;
    
    add_reg_add_reg_2_1 add_reg_5 (.addresult_RNI8MQ7({
        addresult_RNI8MQ7[14]}), .addresult_RNIFE5C({
        \addresult_RNIFE5C[10] }), .signal_data_0_iv_i_2({
        \signal_data_0_iv_i_2[11] , \signal_data_0_iv_i_2[10] , 
        \signal_data_0_iv_i_2[9] , \signal_data_0_iv_i_2[8] , 
        \signal_data_0_iv_i_2[7] , \signal_data_0_iv_i_2[6] , 
        \signal_data_0_iv_i_2[5] , \signal_data_0_iv_i_2[4] }), 
        .addresult_RNIBOIB({\addresult_RNIBOIB[5] }), 
        .signal_data_0_iv_i_5({\signal_data_0_iv_i_5[11] , 
        \signal_data_0_iv_i_5[10] , \signal_data_0_iv_i_5[9] , 
        \signal_data_0_iv_i_5[8] , \signal_data_0_iv_i_5[7] , 
        \signal_data_0_iv_i_5[6] , \signal_data_0_iv_i_5[5] , 
        \signal_data_0_iv_i_5[4] }), .signal_data_iv_0_0_3({
        \signal_data_iv_0_0_3[1] }), .signal_data_iv_0_0_9({
        \signal_data_iv_0_0_9[1] }), .signal_data_iv_0_3_0(
        \signal_data_iv_0_3[0] ), .signal_data_iv_0_3_3(
        \signal_data_iv_0_3[3] ), .signal_data_iv_0_3_2(
        \signal_data_iv_0_3[2] ), .signal_data_iv_0_9_0(
        \signal_data_iv_0_9[0] ), .signal_data_iv_0_9_3(
        \signal_data_iv_0_9[3] ), .signal_data_iv_0_9_2(
        \signal_data_iv_0_9[2] ), .un1_n_s_change_0_1({
        un1_n_s_change_0_1[4], un1_n_s_change_0_1[3], 
        un1_n_s_change_0_1[2], un1_n_s_change_0_1[1], 
        un1_n_s_change_0_1[0]}), .un1_ten_choice_one_0_5({
        \un1_ten_choice_one_0_5[11] , \un1_ten_choice_one_0_5[10] , 
        \un1_ten_choice_one_0_5[9] , \un1_ten_choice_one_0_5[8] , 
        \un1_ten_choice_one_0_5[7] , \un1_ten_choice_one_0_5[6] , 
        \un1_ten_choice_one_0_5[5] , \un1_ten_choice_one_0_5[4] , 
        \un1_ten_choice_one_0_5[3] , \un1_ten_choice_one_0_5[2] , 
        \un1_ten_choice_one_0_5[1] , \un1_ten_choice_one_0_5[0] }), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add), .N_216(
        N_216), .N_249(N_249), .N_184(N_184), .N_200(N_200), .N_255(
        N_255), .N_249_0(N_249_0), .N_233(N_233), .N_262(N_262), 
        .N_111(N_111), .N_95(N_95), .N_250(N_250), .N_87(N_87), .N_210(
        N_210), .N_214(N_214), .N_186(N_186), .N_174(N_174), .N_158(
        N_158), .N_134(N_134), .N_126(N_126), .N_118(N_118), .N_150(
        N_150), .N_235(N_235), .N_202(N_202), .N_218(N_218), .N_223(
        N_223));
    add_reg_add_reg_2_4 add_reg_0 (.un1_n_s_change_0_1({
        un1_n_s_change_0_1[2], un1_n_s_change_0_1[1], 
        un1_n_s_change_0_1[0]}), .signal_data_0_iv_i_5({
        \signal_data_0_iv_i_5[11] , \signal_data_0_iv_i_5[10] , 
        \signal_data_0_iv_i_5[9] , \signal_data_0_iv_i_5[8] , 
        \signal_data_0_iv_i_5[7] , \signal_data_0_iv_i_5[6] , 
        \signal_data_0_iv_i_5[5] , \signal_data_0_iv_i_5[4] }), 
        .signal_data_0_iv_i_3({\signal_data_0_iv_i_3[11] , 
        \signal_data_0_iv_i_3[10] , \signal_data_0_iv_i_3[9] , 
        \signal_data_0_iv_i_3[8] , \signal_data_0_iv_i_3[7] , 
        \signal_data_0_iv_i_3[6] , \signal_data_0_iv_i_3[5] , 
        \signal_data_0_iv_i_3[4] }), .signal_data_0_iv_i_0({
        \signal_data_0_iv_i_0[11] , \signal_data_0_iv_i_0[10] , 
        \signal_data_0_iv_i_0[9] , \signal_data_0_iv_i_0[8] , 
        \signal_data_0_iv_i_0[7] , \signal_data_0_iv_i_0[6] , 
        \signal_data_0_iv_i_0[5] , \signal_data_0_iv_i_0[4] }), 
        .signal_data_iv_0_0_10({\signal_data_iv_0_0_10[1] }), 
        .signal_data_iv_0_0_6({\signal_data_iv_0_0_6[1] }), 
        .signal_data_iv_0_0_13({\signal_data_iv_0_0_13[1] }), 
        .signal_data_iv_0_10_0(\signal_data_iv_0_10[0] ), 
        .signal_data_iv_0_10_3(\signal_data_iv_0_10[3] ), 
        .signal_data_iv_0_10_2(\signal_data_iv_0_10[2] ), 
        .signal_data_iv_0_6_0(\signal_data_iv_0_6[0] ), 
        .signal_data_iv_0_6_3(\signal_data_iv_0_6[3] ), 
        .signal_data_iv_0_6_2(\signal_data_iv_0_6[2] ), 
        .signal_data_iv_0_13_0(\signal_data_iv_0_13[0] ), 
        .signal_data_iv_0_13_3(\signal_data_iv_0_13[3] ), 
        .signal_data_iv_0_13_2(\signal_data_iv_0_13[2] ), 
        .un1_ten_choice_one_0({\un1_ten_choice_one_0[11] , 
        \un1_ten_choice_one_0[10] , \un1_ten_choice_one_0[9] , 
        \un1_ten_choice_one_0[8] , \un1_ten_choice_one_0[7] , 
        \un1_ten_choice_one_0[6] , \un1_ten_choice_one_0[5] , 
        \un1_ten_choice_one_0[4] , \un1_ten_choice_one_0[3] , 
        \un1_ten_choice_one_0[2] , \un1_ten_choice_one_0[1] , 
        \un1_ten_choice_one_0[0] }), .addresult_4_10(addresult_4_2), 
        .addresult_4_8(addresult_4_0), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .signalclkctrl_0_clk_add(
        signalclkctrl_0_clk_add), .N_226(N_226), .N_249(N_249), .N_194(
        N_194), .N_210(N_210_0), .N_254(N_254), .N_249_0(N_249_0), 
        .N_243(N_243), .N_108(N_108), .N_92(N_92), .N_222(N_222), 
        .N_25_i_0(N_25_i_0), .N_20_i_0(N_20_i_0), .N_12_i_0(N_12_i_0), 
        .N_14_i_0(N_14_i_0), .N_16_i_0(N_16_i_0), .N_18_i_0(N_18_i_0), 
        .N_22_i_0(N_22_i_0), .N_27_i_0(N_27_i_0), .N_196(N_196), .N_39(
        N_39), .N_245(N_245), .N_212(N_212), .N_228(N_228), .N_271(
        N_271));
    OR3B \signal_data_0_iv_i_a2_1[12]  (.A(s_addchoice[2]), .B(
        s_addchoice[1]), .C(s_addchoice[3]), .Y(N_252));
    ten_choice_one ten_choice_one_0 (.un1_ten_choice_one_0_7_0(
        \un1_ten_choice_one_0_7[0] ), .un1_ten_choice_one_0_7_2(
        \un1_ten_choice_one_0_7[2] ), .un1_ten_choice_one_0_7_11(
        \un1_ten_choice_one_0_7[11] ), .un1_ten_choice_one_0_7_10(
        \un1_ten_choice_one_0_7[10] ), .un1_ten_choice_one_0_7_9(
        \un1_ten_choice_one_0_7[9] ), .un1_ten_choice_one_0_7_8(
        \un1_ten_choice_one_0_7[8] ), .un1_ten_choice_one_0_7_7(
        \un1_ten_choice_one_0_7[7] ), .un1_ten_choice_one_0_7_6(
        \un1_ten_choice_one_0_7[6] ), .un1_ten_choice_one_0_7_5(
        \un1_ten_choice_one_0_7[5] ), .un1_ten_choice_one_0_7_3(
        \un1_ten_choice_one_0_7[3] ), .un1_ten_choice_one_0_4_3(
        \un1_ten_choice_one_0_4[3] ), .un1_ten_choice_one_0_4_1(
        \un1_ten_choice_one_0_4[1] ), .un1_ten_choice_one_0_4_0(
        \un1_ten_choice_one_0_4[0] ), .un1_ten_choice_one_0_4_11(
        \un1_ten_choice_one_0_4[11] ), .un1_ten_choice_one_0_4_10(
        \un1_ten_choice_one_0_4[10] ), .un1_ten_choice_one_0_4_9(
        \un1_ten_choice_one_0_4[9] ), .un1_ten_choice_one_0_4_8(
        \un1_ten_choice_one_0_4[8] ), .un1_ten_choice_one_0_4_7(
        \un1_ten_choice_one_0_4[7] ), .un1_ten_choice_one_0_4_6(
        \un1_ten_choice_one_0_4[6] ), .un1_ten_choice_one_0_4_5(
        \un1_ten_choice_one_0_4[5] ), .un1_ten_choice_one_0_4_4(
        \un1_ten_choice_one_0_4[4] ), .un1_ten_choice_one_0_3_1(
        \un1_ten_choice_one_0_3[1] ), .un1_ten_choice_one_0_3_0(
        \un1_ten_choice_one_0_3[0] ), .un1_ten_choice_one_0_3_10(
        \un1_ten_choice_one_0_3[10] ), .un1_ten_choice_one_0_3_11(
        \un1_ten_choice_one_0_3[11] ), .un1_ten_choice_one_0_3_9(
        \un1_ten_choice_one_0_3[9] ), .un1_ten_choice_one_0_3_8(
        \un1_ten_choice_one_0_3[8] ), .un1_ten_choice_one_0_3_7(
        \un1_ten_choice_one_0_3[7] ), .un1_ten_choice_one_0_3_6(
        \un1_ten_choice_one_0_3[6] ), .un1_ten_choice_one_0_3_5(
        \un1_ten_choice_one_0_3[5] ), .un1_ten_choice_one_0_3_4(
        \un1_ten_choice_one_0_3[4] ), .un1_ten_choice_one_0_3_3(
        \un1_ten_choice_one_0_3[3] ), .un1_ten_choice_one_0({
        \un1_ten_choice_one_0[11] , \un1_ten_choice_one_0[10] , 
        \un1_ten_choice_one_0[9] , \un1_ten_choice_one_0[8] , 
        \un1_ten_choice_one_0[7] , \un1_ten_choice_one_0[6] , 
        \un1_ten_choice_one_0[5] , \un1_ten_choice_one_0[4] , 
        \un1_ten_choice_one_0[3] , \un1_ten_choice_one_0[2] , 
        \un1_ten_choice_one_0[1] , \un1_ten_choice_one_0[0] }), 
        .un1_ten_choice_one_0_6({\un1_ten_choice_one_0_6[11] , 
        \un1_ten_choice_one_0_6[10] , \un1_ten_choice_one_0_6[9] , 
        \un1_ten_choice_one_0_6[8] , \un1_ten_choice_one_0_6[7] , 
        \un1_ten_choice_one_0_6[6] , \un1_ten_choice_one_0_6[5] , 
        \un1_ten_choice_one_0_6[4] , \un1_ten_choice_one_0_6[3] , 
        \un1_ten_choice_one_0_6[2] , \un1_ten_choice_one_0_6[1] }), 
        .un1_ten_choice_one_0_5({\un1_ten_choice_one_0_5[11] , 
        \un1_ten_choice_one_0_5[10] , \un1_ten_choice_one_0_5[9] , 
        \un1_ten_choice_one_0_5[8] , \un1_ten_choice_one_0_5[7] , 
        \un1_ten_choice_one_0_5[6] , \un1_ten_choice_one_0_5[5] , 
        \un1_ten_choice_one_0_5[4] , \un1_ten_choice_one_0_5[3] , 
        \un1_ten_choice_one_0_5[2] , \un1_ten_choice_one_0_5[1] , 
        \un1_ten_choice_one_0_5[0] }), .un1_ten_choice_one_0_1_2(
        \un1_ten_choice_one_0_1[2] ), .un1_ten_choice_one_0_1_1(
        \un1_ten_choice_one_0_1[1] ), .un1_ten_choice_one_0_1_0(
        \un1_ten_choice_one_0_1[0] ), .un1_ten_choice_one_0_1_8(
        \un1_ten_choice_one_0_1[8] ), .un1_ten_choice_one_0_1_10(
        \un1_ten_choice_one_0_1[10] ), .un1_ten_choice_one_0_1_11(
        \un1_ten_choice_one_0_1[11] ), .un1_ten_choice_one_0_1_9(
        \un1_ten_choice_one_0_1[9] ), .un1_ten_choice_one_0_1_7(
        \un1_ten_choice_one_0_1[7] ), .un1_ten_choice_one_0_1_6(
        \un1_ten_choice_one_0_1[6] ), .un1_ten_choice_one_0_1_5(
        \un1_ten_choice_one_0_1[5] ), .un1_ten_choice_one_0_1_4(
        \un1_ten_choice_one_0_1[4] ), .addrout({\addrout[3] , 
        \addrout[2] , \addrout[1] , \addrout[0] }), 
        .dataeight_0_a2_0_0({\dataeight_0_a2_0_0[0] }), 
        .un1_n_s_change_0_1({un1_n_s_change_0_1[11], 
        un1_n_s_change_0_1[10], un1_n_s_change_0_1[9], 
        un1_n_s_change_0_1[8], un1_n_s_change_0_1[7], 
        un1_n_s_change_0_1[6], un1_n_s_change_0_1[5], 
        un1_n_s_change_0_1[4], un1_n_s_change_0_1[3], 
        un1_n_s_change_0_1[2], un1_n_s_change_0_1[1], 
        un1_n_s_change_0_1[0]}), .un1_ten_choice_one_0_2_0(
        \un1_ten_choice_one_0_2[1] ), .un1_ten_choice_one_0_2_10(
        \un1_ten_choice_one_0_2[11] ), .un1_ten_choice_one_0_2_9(
        \un1_ten_choice_one_0_2[10] ), .un1_ten_choice_one_0_2_8(
        \un1_ten_choice_one_0_2[9] ), .un1_ten_choice_one_0_2_7(
        \un1_ten_choice_one_0_2[8] ), .un1_ten_choice_one_0_2_6(
        \un1_ten_choice_one_0_2[7] ), .un1_ten_choice_one_0_2_5(
        \un1_ten_choice_one_0_2[6] ), .un1_ten_choice_one_0_2_4(
        \un1_ten_choice_one_0_2[5] ), .un1_ten_choice_one_0_2_3(
        \un1_ten_choice_one_0_2[4] ), .un1_ten_choice_one_0_2_2(
        \un1_ten_choice_one_0_2[3] ), .N_214(N_214), .N_212(N_212_0), 
        .N_211(N_211), .N_217(N_217), .N_219(N_219), .N_222(N_222), 
        .N_221(N_221_0), .N_223(N_223), .N_224(N_224_0), .N_216(
        N_216_0), .N_213(N_213), .N_220(N_220_0), .N_210(N_210), 
        .N_215(N_215));
    add_reg_add_reg_2_7 add_reg_4 (.addresult_RNIVJME({
        \addresult_RNIVJME[4] }), .signal_data_0_iv_i_2({
        \signal_data_0_iv_i_2[11] , \signal_data_0_iv_i_2[10] , 
        \signal_data_0_iv_i_2[9] , \signal_data_0_iv_i_2[8] , 
        \signal_data_0_iv_i_2[7] , \signal_data_0_iv_i_2[6] , 
        \signal_data_0_iv_i_2[5] , \signal_data_0_iv_i_2[4] }), 
        .signal_data_iv_0_0_3({\signal_data_iv_0_0_3[1] }), 
        .signal_data_iv_0_3_0(\signal_data_iv_0_3[0] ), 
        .signal_data_iv_0_3_3(\signal_data_iv_0_3[3] ), 
        .signal_data_iv_0_3_2(\signal_data_iv_0_3[2] ), .ADC_c({
        ADC_c[2], ADC_c[1], ADC_c[0]}), .un1_n_s_change_0_1({
        un1_n_s_change_0_1[3], un1_n_s_change_0_1[2]}), 
        .un1_ten_choice_one_0_4_0(\un1_ten_choice_one_0_4[0] ), 
        .un1_ten_choice_one_0_4_3(\un1_ten_choice_one_0_4[3] ), 
        .un1_ten_choice_one_0_4_1(\un1_ten_choice_one_0_4[1] ), 
        .un1_ten_choice_one_0_4_4(\un1_ten_choice_one_0_4[4] ), 
        .un1_ten_choice_one_0_4_5(\un1_ten_choice_one_0_4[5] ), 
        .un1_ten_choice_one_0_4_7(\un1_ten_choice_one_0_4[7] ), 
        .un1_ten_choice_one_0_4_8(\un1_ten_choice_one_0_4[8] ), 
        .un1_ten_choice_one_0_4_9(\un1_ten_choice_one_0_4[9] ), 
        .un1_ten_choice_one_0_4_10(\un1_ten_choice_one_0_4[10] ), 
        .un1_ten_choice_one_0_4_11(\un1_ten_choice_one_0_4[11] ), 
        .un1_ten_choice_one_0_4_6(\un1_ten_choice_one_0_4[6] ), 
        .un1_add_reg_4_i_2(un1_add_reg_4_i_2), .un1_add_reg_4_i_0(
        un1_add_reg_4_i_0), .s_acq_change_0_s_rst(s_acq_change_0_s_rst)
        , .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add), .N_218(
        N_218), .N_186(N_186), .N_88(N_88), .N_104(N_104), .N_249(
        N_249), .N_202(N_202), .N_250(N_250), .N_249_0(N_249_0), 
        .N_235(N_235), .N_212(N_212_0), .N_211(N_211), .N_188(N_188), 
        .N_177(N_177), .N_145(N_145), .N_137(N_137), .N_129(N_129), 
        .N_121(N_121), .N_153(N_153), .N_169(N_169), .N_253(N_253), 
        .N_237(N_237), .N_204(N_204), .N_220(N_220), .N_263(N_263), 
        .top_code_0_n_s_ctrl_0(top_code_0_n_s_ctrl_0), .N_217(N_217));
    s_clk_div4 s_clk_div4_0 (.s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .ddsclkout_c(ddsclkout_c), .clkout(
        clkout), .scan_scale_sw_0_s_start(scan_scale_sw_0_s_start), 
        .signalclkctrl_0_entop(signalclkctrl_0_entop));
    NOR2 \signal_data_iv_0_a2_3[0]  (.A(N_253), .B(N_33), .Y(N_263));
    OR2A \signal_data_0_iv_i_o17[12]  (.A(s_addchoice[0]), .B(
        s_addchoice[4]), .Y(N_33));
    OR3A \signal_data_0_iv_i_a2_2[12]  (.A(s_addchoice[3]), .B(
        s_addchoice[2]), .C(s_addchoice[1]), .Y(N_253));
    OR3B \signal_data_0_iv_i_a2_4[12]  (.A(s_addchoice[2]), .B(
        s_addchoice[3]), .C(s_addchoice[1]), .Y(N_255));
    VCC VCC_i (.Y(VCC));
    ctrl_addr ctrl_addr_0 (.s_periodnum({s_periodnum[3], 
        s_periodnum[2], s_periodnum[1], s_periodnum[0]}), .addrout({
        \addrout[3] , \addrout[2] , \addrout[1] , \addrout[0] }), 
        .s_acq_change_0_s_load_0(s_acq_change_0_s_load_0), .GLA(GLA), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add));
    OR3 G_1_0_o2 (.A(s_addchoice[2]), .B(s_addchoice[3]), .C(
        s_addchoice[1]), .Y(N_39));
    OR3C \signal_data_0_iv_i_a2_5[12]  (.A(s_addchoice[2]), .B(
        s_addchoice[3]), .C(s_addchoice[1]), .Y(N_256));
    NOR2 \signal_data_iv_0_a2_7[0]  (.A(N_256), .B(N_33), .Y(N_267));
    NOR2 \signal_data_iv_0_a2_6[0]  (.A(N_252), .B(N_33), .Y(N_266));
    OR3A \signal_data_0_iv_i_a2_0[12]  (.A(s_addchoice[2]), .B(
        s_addchoice[3]), .C(s_addchoice[1]), .Y(N_251));
    OR3A \signal_data_0_iv_i_a2_3[12]  (.A(s_addchoice[1]), .B(
        s_addchoice[2]), .C(s_addchoice[3]), .Y(N_254));
    OR2 \signal_data_iv_0_a2_14[0]  (.A(s_addchoice[4]), .B(
        s_addchoice[0]), .Y(N_249));
    NOR2 \signal_data_iv_0_a2[0]  (.A(N_251), .B(N_33), .Y(N_259));
    GND GND_i (.Y(GND));
    OR2 \signal_data_iv_0_a2_14_0[0]  (.A(s_addchoice[4]), .B(
        s_addchoice[0]), .Y(N_249_0));
    add_reg_add_reg_2_3 add_reg_1 (.addresult_RNIDU3E({
        \addresult_RNIDU3E[4] }), .signal_data_iv_0_0_6({
        \signal_data_iv_0_0_6[1] }), .signal_data_iv_0_6_0(
        \signal_data_iv_0_6[0] ), .signal_data_iv_0_6_3(
        \signal_data_iv_0_6[3] ), .signal_data_iv_0_6_2(
        \signal_data_iv_0_6[2] ), .un1_n_s_change_0_1({
        un1_n_s_change_0_1[3], un1_n_s_change_0_1[2], 
        un1_n_s_change_0_1[1], un1_n_s_change_0_1[0]}), 
        .un1_ten_choice_one_0_1_0(\un1_ten_choice_one_0_1[0] ), 
        .un1_ten_choice_one_0_1_2(\un1_ten_choice_one_0_1[2] ), 
        .un1_ten_choice_one_0_1_10(\un1_ten_choice_one_0_1[10] ), 
        .un1_ten_choice_one_0_1_5(\un1_ten_choice_one_0_1[5] ), 
        .un1_ten_choice_one_0_1_9(\un1_ten_choice_one_0_1[9] ), 
        .un1_ten_choice_one_0_1_7(\un1_ten_choice_one_0_1[7] ), 
        .un1_ten_choice_one_0_1_1(\un1_ten_choice_one_0_1[1] ), 
        .un1_ten_choice_one_0_1_8(\un1_ten_choice_one_0_1[8] ), 
        .un1_ten_choice_one_0_1_4(\un1_ten_choice_one_0_1[4] ), 
        .un1_ten_choice_one_0_1_6(\un1_ten_choice_one_0_1[6] ), 
        .un1_ten_choice_one_0_1_11(\un1_ten_choice_one_0_1[11] ), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add), .N_249(
        N_249), .N_224(N_224), .N_91(N_91), .N_107(N_107), .N_192(
        N_192), .N_208(N_208), .N_251(N_251), .N_249_0(N_249_0), 
        .N_241(N_241), .N_179(N_179), .N_171(N_171), .N_155(N_155), 
        .N_147(N_147), .N_139(N_139), .N_131(N_131), .N_123(N_123), 
        .N_115(N_115), .N_254(N_254), .N_99(N_99), .N_194(N_194), 
        .N_243(N_243), .N_210_0(N_210_0), .N_226(N_226), .N_273(N_273), 
        .N_213(N_213), .N_210(N_210), .N_216(N_216_0));
    AX1B G_1_0 (.A(N_39), .B(s_addchoice[0]), .C(s_addchoice[4]), .Y(
        \signal_data_en[9] ));
    NOR2A G_1_0_a2_0 (.A(s_addchoice[4]), .B(N_39), .Y(
        G_1_0_a2_0_net_1));
    NOR2 \signal_data_iv_0_a2_10[0]  (.A(N_255), .B(N_33), .Y(N_270));
    add_reg_add_reg_2_6 add_reg_6 (.addresult_RNIJE5C({
        addresult_RNIJE5C[14]}), .addresult_RNIFE5C({
        \addresult_RNIFE5C[10] }), .addresult_RNIBOIB({
        \addresult_RNIBOIB[5] }), .addresult_0_15(addresult_0_2), 
        .addresult_0_13(addresult_0_0), .signal_data_iv_0_0_1({
        \signal_data_iv_0_0_1[1] }), .signal_data_iv_0_1_0(
        \signal_data_iv_0_1[0] ), .signal_data_iv_0_1_3(
        \signal_data_iv_0_1[3] ), .signal_data_iv_0_1_2(
        \signal_data_iv_0_1[2] ), .un1_n_s_change_0_1({
        un1_n_s_change_0_1[2], un1_n_s_change_0_1[1], 
        un1_n_s_change_0_1[0]}), .un1_ten_choice_one_0_6({
        \un1_ten_choice_one_0_6[11] , \un1_ten_choice_one_0_6[10] , 
        \un1_ten_choice_one_0_6[9] , \un1_ten_choice_one_0_6[8] , 
        \un1_ten_choice_one_0_6[7] , \un1_ten_choice_one_0_6[6] , 
        \un1_ten_choice_one_0_6[5] , \un1_ten_choice_one_0_6[4] , 
        \un1_ten_choice_one_0_6[3] , \un1_ten_choice_one_0_6[2] , 
        \un1_ten_choice_one_0_6[1] }), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .signalclkctrl_0_clk_add(
        signalclkctrl_0_clk_add), .N_214(N_214_0), .N_182(N_182), 
        .N_221(N_221_0), .N_249(N_249), .N_198(N_198), .N_256(N_256), 
        .N_249_0(N_249_0), .N_231(N_231), .N_174(N_174), .N_158(N_158), 
        .N_150(N_150), .N_134(N_134), .N_126(N_126), .N_118(N_118), 
        .N_255(N_255), .N_86(N_86), .N_210(N_210), .N_212(N_212_0), 
        .N_184(N_184), .N_233(N_233), .N_200(N_200), .N_216(N_216), 
        .N_270(N_270));
    add_reg_add_reg_2_5 add_reg_7 (.s_addchoice({s_addchoice[0]}), 
        .signal_data_iv_0_0_13({\signal_data_iv_0_0_13[1] }), 
        .signal_data_en({\signal_data_en[9] }), .signal_data_iv_0_13_2(
        \signal_data_iv_0_13[2] ), .signal_data_iv_0_13_3(
        \signal_data_iv_0_13[3] ), .signal_data_iv_0_13_0(
        \signal_data_iv_0_13[0] ), .un1_signal_acq_0({
        un1_signal_acq_0[3], un1_signal_acq_0[2], un1_signal_acq_0[1], 
        un1_signal_acq_0[0]}), .dataeight_0_a2_0_0({
        \dataeight_0_a2_0_0[0] }), .signal_data_0_iv_i_0({
        \signal_data_0_iv_i_0[11] , \signal_data_0_iv_i_0[10] , 
        \signal_data_0_iv_i_0[9] , \signal_data_0_iv_i_0[8] , 
        \signal_data_0_iv_i_0[7] , \signal_data_0_iv_i_0[6] , 
        \signal_data_0_iv_i_0[5] , \signal_data_0_iv_i_0[4] }), 
        .signal_data_iv_0_0_9({\signal_data_iv_0_0_9[1] }), 
        .signal_data_iv_0_0_1({\signal_data_iv_0_0_1[1] }), 
        .signal_data_iv_0_9_0(\signal_data_iv_0_9[0] ), 
        .signal_data_iv_0_9_3(\signal_data_iv_0_9[3] ), 
        .signal_data_iv_0_9_2(\signal_data_iv_0_9[2] ), 
        .signal_data_iv_0_1_0(\signal_data_iv_0_1[0] ), 
        .signal_data_iv_0_1_3(\signal_data_iv_0_1[3] ), 
        .signal_data_iv_0_1_2(\signal_data_iv_0_1[2] ), .addresult_14(
        addresult[14]), .addresult_13(addresult[13]), .addresult_15(
        addresult[15]), .addresult_12(addresult[12]), 
        .un1_ten_choice_one_0_7_2(\un1_ten_choice_one_0_7[2] ), 
        .un1_ten_choice_one_0_7_3(\un1_ten_choice_one_0_7[3] ), 
        .un1_ten_choice_one_0_7_5(\un1_ten_choice_one_0_7[5] ), 
        .un1_ten_choice_one_0_7_6(\un1_ten_choice_one_0_7[6] ), 
        .un1_ten_choice_one_0_7_7(\un1_ten_choice_one_0_7[7] ), 
        .un1_ten_choice_one_0_7_8(\un1_ten_choice_one_0_7[8] ), 
        .un1_ten_choice_one_0_7_9(\un1_ten_choice_one_0_7[9] ), 
        .un1_ten_choice_one_0_7_10(\un1_ten_choice_one_0_7[10] ), 
        .un1_ten_choice_one_0_7_11(\un1_ten_choice_one_0_7[11] ), 
        .un1_ten_choice_one_0_7_0(\un1_ten_choice_one_0_7[0] ), 
        .un1_n_s_change_0_1({un1_n_s_change_0_1[4], 
        un1_n_s_change_0_1[3], un1_n_s_change_0_1[2], 
        un1_n_s_change_0_1[1], un1_n_s_change_0_1[0]}), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add), .N_228(
        N_228), .N_245(N_245), .N_196(N_196), .G_1_0_a2_0(
        G_1_0_a2_0_net_1), .N_212(N_212), .N_213(N_213), .N_182(N_182), 
        .N_33(N_33), .N_256(N_256), .N_231(N_231), .N_198(N_198), 
        .N_214(N_214_0), .N_267(N_267), .N_220(N_220_0));
    NOR2 \signal_data_iv_0_a2_2[0]  (.A(N_250), .B(N_33), .Y(N_262));
    NOR2 \signal_data_iv_0_a2_11[0]  (.A(N_39), .B(N_33), .Y(N_271));
    add_reg_add_reg_2 add_reg_2 (.addresult_RNI5DQA({
        addresult_RNI5DQA[12]}), .addresult_RNI7DQA({
        addresult_RNI7DQA[14]}), .addresult_5_10(addresult_5_2), 
        .addresult_5_8(addresult_5_0), .addresult_RNIDU3E({
        \addresult_RNIDU3E[4] }), .signal_data_0_iv_i_3({
        \signal_data_0_iv_i_3[11] , \signal_data_0_iv_i_3[10] , 
        \signal_data_0_iv_i_3[9] , \signal_data_0_iv_i_3[8] , 
        \signal_data_0_iv_i_3[7] , \signal_data_0_iv_i_3[6] , 
        \signal_data_0_iv_i_3[5] , \signal_data_0_iv_i_3[4] }), 
        .signal_data_iv_0_0_10({\signal_data_iv_0_0_10[1] }), 
        .signal_data_iv_0_10_0(\signal_data_iv_0_10[0] ), 
        .signal_data_iv_0_10_3(\signal_data_iv_0_10[3] ), 
        .signal_data_iv_0_10_2(\signal_data_iv_0_10[2] ), 
        .un1_ten_choice_one_0_2_0(\un1_ten_choice_one_0_2[1] ), 
        .un1_ten_choice_one_0_2_2(\un1_ten_choice_one_0_2[3] ), 
        .un1_ten_choice_one_0_2_3(\un1_ten_choice_one_0_2[4] ), 
        .un1_ten_choice_one_0_2_4(\un1_ten_choice_one_0_2[5] ), 
        .un1_ten_choice_one_0_2_5(\un1_ten_choice_one_0_2[6] ), 
        .un1_ten_choice_one_0_2_7(\un1_ten_choice_one_0_2[8] ), 
        .un1_ten_choice_one_0_2_8(\un1_ten_choice_one_0_2[9] ), 
        .un1_ten_choice_one_0_2_9(\un1_ten_choice_one_0_2[10] ), 
        .un1_ten_choice_one_0_2_10(\un1_ten_choice_one_0_2[11] ), 
        .un1_ten_choice_one_0_2_6(\un1_ten_choice_one_0_2[7] ), 
        .un1_n_s_change_0_1({un1_n_s_change_0_1[2], 
        un1_n_s_change_0_1[1], un1_n_s_change_0_1[0]}), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add), .N_249(
        N_249), .N_252(N_252), .N_249_0(N_249_0), .N_215(N_215), 
        .N_210(N_210), .N_192(N_192), .N_189(N_189), .N_179(N_179), 
        .N_147(N_147), .N_139(N_139), .N_131(N_131), .N_123(N_123), 
        .N_155(N_155), .N_171(N_171), .N_251(N_251), .N_241(N_241), 
        .N_238(N_238), .N_208(N_208), .N_205(N_205), .N_224_0(N_224), 
        .N_259(N_259), .N_221(N_221), .N_224(N_224_0));
    OR3B \signal_data_0_iv_i_a2[12]  (.A(s_addchoice[3]), .B(
        s_addchoice[1]), .C(s_addchoice[2]), .Y(N_250));
    add_reg_add_reg_2_2 add_reg_3 (.addresult_RNIVJME({
        \addresult_RNIVJME[4] }), .un1_n_s_change_0_1({
        un1_n_s_change_0_1[2], un1_n_s_change_0_1[1], 
        un1_n_s_change_0_1[0]}), .un1_ten_choice_one_0_3_0(
        \un1_ten_choice_one_0_3[0] ), .un1_ten_choice_one_0_3_1(
        \un1_ten_choice_one_0_3[1] ), .un1_ten_choice_one_0_3_3(
        \un1_ten_choice_one_0_3[3] ), .un1_ten_choice_one_0_3_10(
        \un1_ten_choice_one_0_3[10] ), .un1_ten_choice_one_0_3_4(
        \un1_ten_choice_one_0_3[4] ), .un1_ten_choice_one_0_3_6(
        \un1_ten_choice_one_0_3[6] ), .un1_ten_choice_one_0_3_7(
        \un1_ten_choice_one_0_3[7] ), .un1_ten_choice_one_0_3_8(
        \un1_ten_choice_one_0_3[8] ), .un1_ten_choice_one_0_3_9(
        \un1_ten_choice_one_0_3[9] ), .un1_ten_choice_one_0_3_11(
        \un1_ten_choice_one_0_3[11] ), .un1_ten_choice_one_0_3_5(
        \un1_ten_choice_one_0_3[5] ), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .signalclkctrl_0_clk_add(
        signalclkctrl_0_clk_add), .N_249(N_249), .N_220(N_220), .N_221(
        N_221), .N_205(N_205), .N_89(N_89), .N_105(N_105), .N_204(
        N_204), .N_189(N_189), .N_266(N_266), .N_238(N_238), .N_237(
        N_237), .N_253(N_253), .N_249_0(N_249_0), .N_188(N_188), 
        .N_177(N_177), .N_169(N_169), .N_153(N_153), .N_145(N_145), 
        .N_137(N_137), .N_129(N_129), .N_121(N_121), .N_113(N_113), 
        .N_252(N_252), .N_97(N_97), .N_219(N_219));
    NOR2 \signal_data_iv_0_a2_13[0]  (.A(N_254), .B(N_33), .Y(N_273));
    signalclkctrl signalclkctrl_0 (.s_acqnum({s_acqnum[15], 
        s_acqnum[14], s_acqnum[13], s_acqnum[12], s_acqnum[11], 
        s_acqnum[10], s_acqnum[9], s_acqnum[8], s_acqnum[7], 
        s_acqnum[6], s_acqnum[5], s_acqnum[4], s_acqnum[3], 
        s_acqnum[2], s_acqnum[1], s_acqnum[0]}), .s_periodnum({
        s_periodnum[3], s_periodnum[2], s_periodnum[1], s_periodnum[0]})
        , .s_stripnum({s_stripnum[11], s_stripnum[10], s_stripnum[9], 
        s_stripnum[8], s_stripnum[7], s_stripnum[6], s_stripnum[5], 
        s_stripnum[4], s_stripnum[3], s_stripnum[2], s_stripnum[1], 
        s_stripnum[0]}), .s_acq_change_0_s_load_0(
        s_acq_change_0_s_load_0), .s_acq_change_0_s_load(
        s_acq_change_0_s_load), .GLA(GLA), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .signalclkctrl_0_entop(
        signalclkctrl_0_entop), .signal_acq_0_Signal_acq_clk(
        signal_acq_0_Signal_acq_clk), .clkout(clkout), 
        .signalclkctrl_0_clk_add(signalclkctrl_0_clk_add));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module n_s_change(
       un1_signal_acq_0,
       dataout_0_2,
       dataout_0_3,
       dataout_0_1,
       dataout_0_5,
       dataout_0_11,
       dataout_0_7,
       dataout_0_8,
       dataout_0_6,
       dataout_0_0_d0,
       dataout_0_10,
       dataout_0_9,
       dataout_0_4,
       dataout_0_0,
       addresult_RNI5DQA,
       addresult_RNIJE5C,
       addresult_RNI8MQ7,
       addresult_RNI7DQA,
       addresult,
       addresult_0_0,
       addresult_0_2,
       un1_add_reg_4_i_0,
       un1_add_reg_4_i_2,
       addresult_5_0,
       addresult_5_2,
       addresult_4_0,
       addresult_4_2,
       MX2_RD_2_inst,
       MX2_RD_3_inst,
       MX2_RD_1_inst,
       MX2_RD_5_inst,
       N_25_i_0,
       top_code_0_n_s_ctrl,
       MX2_RD_11_inst,
       N_20_i_0,
       MX2_RD_7_inst,
       N_12_i_0,
       s_clk_div4_0_clkout,
       signal_acq_0_Signal_acq_clk,
       Signal_Noise_Acq_0_acq_clk,
       top_code_0_n_s_ctrl_1,
       MX2_RD_8_inst,
       N_14_i_0,
       MX2_RD_6_inst,
       N_27_i_0,
       MX2_RD_0_inst,
       MX2_RD_10_inst,
       N_18_i_0,
       MX2_RD_9_inst,
       N_16_i_0,
       MX2_RD_4_inst,
       N_22_i_0,
       N_89,
       N_88,
       N_92,
       N_86,
       N_87,
       N_91,
       N_95,
       N_97,
       N_99,
       N_105,
       N_104,
       N_108,
       N_107,
       N_33,
       N_256,
       N_111,
       N_255,
       N_113,
       N_253,
       N_115,
       N_251,
       top_code_0_n_s_ctrl_0,
       N_39
    );
input  [3:0] un1_signal_acq_0;
output dataout_0_2;
output dataout_0_3;
output dataout_0_1;
output dataout_0_5;
output dataout_0_11;
output dataout_0_7;
output dataout_0_8;
output dataout_0_6;
output dataout_0_0_d0;
output dataout_0_10;
output dataout_0_9;
output dataout_0_4;
output [15:12] dataout_0_0;
input  [12:12] addresult_RNI5DQA;
input  [14:14] addresult_RNIJE5C;
input  [14:14] addresult_RNI8MQ7;
input  [14:14] addresult_RNI7DQA;
input  [15:12] addresult;
input  addresult_0_0;
input  addresult_0_2;
input  un1_add_reg_4_i_0;
input  un1_add_reg_4_i_2;
input  addresult_5_0;
input  addresult_5_2;
input  addresult_4_0;
input  addresult_4_2;
input  MX2_RD_2_inst;
input  MX2_RD_3_inst;
input  MX2_RD_1_inst;
input  MX2_RD_5_inst;
input  N_25_i_0;
input  top_code_0_n_s_ctrl;
input  MX2_RD_11_inst;
input  N_20_i_0;
input  MX2_RD_7_inst;
input  N_12_i_0;
input  s_clk_div4_0_clkout;
input  signal_acq_0_Signal_acq_clk;
output Signal_Noise_Acq_0_acq_clk;
input  top_code_0_n_s_ctrl_1;
input  MX2_RD_8_inst;
input  N_14_i_0;
input  MX2_RD_6_inst;
input  N_27_i_0;
input  MX2_RD_0_inst;
input  MX2_RD_10_inst;
input  N_18_i_0;
input  MX2_RD_9_inst;
input  N_16_i_0;
input  MX2_RD_4_inst;
input  N_22_i_0;
input  N_89;
input  N_88;
input  N_92;
input  N_86;
input  N_87;
input  N_91;
input  N_95;
input  N_97;
input  N_99;
input  N_105;
input  N_104;
input  N_108;
input  N_107;
input  N_33;
input  N_256;
input  N_111;
input  N_255;
input  N_113;
input  N_253;
input  N_115;
input  N_251;
input  top_code_0_n_s_ctrl_0;
input  N_39;

    wire \dataout_7[15]_net_1 , \dataout_1[15]_net_1 , 
        \dataout_0[15]_net_1 , \dataout_4[15]_net_1 , 
        \dataout_3[15]_net_1 , \dataout_2[15]_net_1 , 
        \dataout_6[14]_net_1 , \dataout_2[14]_net_1 , 
        \dataout_5[14]_net_1 , \dataout_0[14]_net_1 , 
        \dataout_4[14]_net_1 , \dataout_7[13]_net_1 , 
        \dataout_1[13]_net_1 , \dataout_0[13]_net_1 , 
        \dataout_4[13]_net_1 , \dataout_3[13]_net_1 , 
        \dataout_2[13]_net_1 , \dataout_6[12]_net_1 , 
        \dataout_2[12]_net_1 , \dataout_5[12]_net_1 , 
        \dataout_0[12]_net_1 , \dataout_4[12]_net_1 , GND, VCC, GND_0, 
        VCC_0;
    
    MX2 \dataout[6]  (.A(N_27_i_0), .B(MX2_RD_6_inst), .S(
        top_code_0_n_s_ctrl_0), .Y(dataout_0_6));
    OA1A \dataout_2[13]  (.A(un1_add_reg_4_i_0), .B(N_253), .C(N_97), 
        .Y(\dataout_2[13]_net_1 ));
    MX2 \dataout[11]  (.A(N_20_i_0), .B(MX2_RD_11_inst), .S(
        top_code_0_n_s_ctrl), .Y(dataout_0_11));
    OA1 \dataout_3[15]  (.A(N_251), .B(addresult_5_2), .C(N_115), .Y(
        \dataout_3[15]_net_1 ));
    MX2 \dataout[1]  (.A(un1_signal_acq_0[1]), .B(MX2_RD_1_inst), .S(
        top_code_0_n_s_ctrl), .Y(dataout_0_1));
    NOR3C \dataout[13]  (.A(\dataout_3[13]_net_1 ), .B(
        \dataout_2[13]_net_1 ), .C(\dataout_7[13]_net_1 ), .Y(
        dataout_0_0[13]));
    NOR3C \dataout_5[14]  (.A(addresult_RNI8MQ7[14]), .B(
        addresult_RNIJE5C[14]), .C(\dataout_0[14]_net_1 ), .Y(
        \dataout_5[14]_net_1 ));
    OA1B \dataout_4[13]  (.A(N_39), .B(addresult_4_0), .C(
        top_code_0_n_s_ctrl_0), .Y(\dataout_4[13]_net_1 ));
    MX2 \dataout[0]  (.A(un1_signal_acq_0[0]), .B(MX2_RD_0_inst), .S(
        top_code_0_n_s_ctrl_0), .Y(dataout_0_0_d0));
    VCC VCC_i (.Y(VCC));
    OA1A \dataout_2[15]  (.A(un1_add_reg_4_i_2), .B(N_253), .C(N_113), 
        .Y(\dataout_2[15]_net_1 ));
    NOR2B \dataout_2[12]  (.A(N_88), .B(N_89), .Y(
        \dataout_2[12]_net_1 ));
    MX2 \dataout[10]  (.A(N_18_i_0), .B(MX2_RD_10_inst), .S(
        top_code_0_n_s_ctrl_0), .Y(dataout_0_10));
    MX2 \dataout[4]  (.A(N_22_i_0), .B(MX2_RD_4_inst), .S(
        top_code_0_n_s_ctrl_0), .Y(dataout_0_4));
    MX2A acq_clk (.A(signal_acq_0_Signal_acq_clk), .B(
        s_clk_div4_0_clkout), .S(top_code_0_n_s_ctrl_1), .Y(
        Signal_Noise_Acq_0_acq_clk));
    NOR3C \dataout[15]  (.A(\dataout_3[15]_net_1 ), .B(
        \dataout_2[15]_net_1 ), .C(\dataout_7[15]_net_1 ), .Y(
        dataout_0_0[15]));
    NOR3C \dataout_7[13]  (.A(\dataout_1[13]_net_1 ), .B(
        \dataout_0[13]_net_1 ), .C(\dataout_4[13]_net_1 ), .Y(
        \dataout_7[13]_net_1 ));
    MX2 \dataout[9]  (.A(N_16_i_0), .B(MX2_RD_9_inst), .S(
        top_code_0_n_s_ctrl_0), .Y(dataout_0_9));
    OA1B \dataout_4[15]  (.A(N_39), .B(addresult_4_2), .C(
        top_code_0_n_s_ctrl_0), .Y(\dataout_4[15]_net_1 ));
    NOR2A \dataout_4[12]  (.A(N_92), .B(top_code_0_n_s_ctrl_0), .Y(
        \dataout_4[12]_net_1 ));
    NOR3C \dataout_6[12]  (.A(N_91), .B(addresult_RNI5DQA[12]), .C(
        \dataout_2[12]_net_1 ), .Y(\dataout_6[12]_net_1 ));
    NOR2B \dataout_2[14]  (.A(N_104), .B(N_105), .Y(
        \dataout_2[14]_net_1 ));
    OA1B \dataout_0[13]  (.A(N_256), .B(addresult[13]), .C(N_33), .Y(
        \dataout_0[13]_net_1 ));
    NOR3C \dataout_7[15]  (.A(\dataout_1[15]_net_1 ), .B(
        \dataout_0[15]_net_1 ), .C(\dataout_4[15]_net_1 ), .Y(
        \dataout_7[15]_net_1 ));
    OA1 \dataout_1[13]  (.A(N_255), .B(addresult_0_0), .C(N_95), .Y(
        \dataout_1[13]_net_1 ));
    GND GND_i (.Y(GND));
    NOR3C \dataout[14]  (.A(\dataout_5[14]_net_1 ), .B(
        \dataout_4[14]_net_1 ), .C(\dataout_6[14]_net_1 ), .Y(
        dataout_0_0[14]));
    NOR2A \dataout_4[14]  (.A(N_108), .B(top_code_0_n_s_ctrl_0), .Y(
        \dataout_4[14]_net_1 ));
    NOR3C \dataout_6[14]  (.A(N_107), .B(addresult_RNI7DQA[14]), .C(
        \dataout_2[14]_net_1 ), .Y(\dataout_6[14]_net_1 ));
    MX2 \dataout[8]  (.A(N_14_i_0), .B(MX2_RD_8_inst), .S(
        top_code_0_n_s_ctrl_1), .Y(dataout_0_8));
    MX2 \dataout[3]  (.A(un1_signal_acq_0[3]), .B(MX2_RD_3_inst), .S(
        top_code_0_n_s_ctrl), .Y(dataout_0_3));
    OA1B \dataout_0[15]  (.A(N_256), .B(addresult[15]), .C(N_33), .Y(
        \dataout_0[15]_net_1 ));
    OA1B \dataout_0[12]  (.A(N_256), .B(addresult[12]), .C(N_33), .Y(
        \dataout_0[12]_net_1 ));
    OA1 \dataout_1[15]  (.A(N_255), .B(addresult_0_2), .C(N_111), .Y(
        \dataout_1[15]_net_1 ));
    MX2 \dataout[7]  (.A(N_12_i_0), .B(MX2_RD_7_inst), .S(
        top_code_0_n_s_ctrl_1), .Y(dataout_0_7));
    NOR3C \dataout[12]  (.A(\dataout_5[12]_net_1 ), .B(
        \dataout_4[12]_net_1 ), .C(\dataout_6[12]_net_1 ), .Y(
        dataout_0_0[12]));
    MX2 \dataout[2]  (.A(un1_signal_acq_0[2]), .B(MX2_RD_2_inst), .S(
        top_code_0_n_s_ctrl), .Y(dataout_0_2));
    MX2 \dataout[5]  (.A(N_25_i_0), .B(MX2_RD_5_inst), .S(
        top_code_0_n_s_ctrl), .Y(dataout_0_5));
    OA1 \dataout_3[13]  (.A(N_251), .B(addresult_5_0), .C(N_99), .Y(
        \dataout_3[13]_net_1 ));
    OA1B \dataout_0[14]  (.A(N_256), .B(addresult[14]), .C(N_33), .Y(
        \dataout_0[14]_net_1 ));
    NOR3C \dataout_5[12]  (.A(N_87), .B(N_86), .C(
        \dataout_0[12]_net_1 ), .Y(\dataout_5[12]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module n_rdclk_syn(
       n_rdclk,
       GLA,
       XRD_c,
       n_acq_change_0_n_rst_n_0,
       top_code_0_n_rd_en
    );
output n_rdclk;
input  GLA;
input  XRD_c;
input  n_acq_change_0_n_rst_n_0;
input  top_code_0_n_rd_en;

    wire n_rdclk_RNO_net_1, un1_clk_wire, clk_reg1_RNO_net_1, 
        clk_reg2_RNO_net_1, clk_reg1_net_1, clk_reg2_net_1, GND, VCC, 
        GND_0, VCC_0;
    
    NOR3B n_rdclk_RNO (.A(top_code_0_n_rd_en), .B(
        n_acq_change_0_n_rst_n_0), .C(un1_clk_wire), .Y(
        n_rdclk_RNO_net_1));
    NOR2B clk_reg2_RNO (.A(n_acq_change_0_n_rst_n_0), .B(
        clk_reg1_net_1), .Y(clk_reg2_RNO_net_1));
    DFN1 n_rdclk_inst_1 (.D(n_rdclk_RNO_net_1), .CLK(GLA), .Q(n_rdclk));
    DFN1 clk_reg2 (.D(clk_reg2_RNO_net_1), .CLK(GLA), .Q(
        clk_reg2_net_1));
    NOR2B clk_reg1_RNO (.A(n_acq_change_0_n_rst_n_0), .B(XRD_c), .Y(
        clk_reg1_RNO_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2A n_rdclk_RNO_0 (.A(clk_reg2_net_1), .B(clk_reg1_net_1), .Y(
        un1_clk_wire));
    DFN1 clk_reg1 (.D(clk_reg1_RNO_net_1), .CLK(GLA), .Q(
        clk_reg1_net_1));
    VCC VCC_i (.Y(VCC));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    
endmodule


module noise_addr_noise_addr_0(
       addr_0,
       n_acq_change_0_n_rst_n,
       n_acq_change_0_n_rst_n_0,
       s_clk_div4_0_clkout
    );
output [11:0] addr_0;
input  n_acq_change_0_n_rst_n;
input  n_acq_change_0_n_rst_n_0;
input  s_clk_div4_0_clkout;

    wire \un1_noise_addr_0_i[0] , addr_n11, addr_c9, addr_n10, addr_n9, 
        addr_c8, addr_n8, addr_c6, addr_n7, addr_n6, addr_c4, addr_n5, 
        addr_n4, addr_c2, addr_n3, addr_n2, addr_n1, GND, VCC, GND_0, 
        VCC_0;
    
    DFN0C0 \addr[6]  (.D(addr_n6), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[6]));
    DFN0C0 \addr[11]  (.D(addr_n11), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[11]));
    XNOR2 \addr_RNO[7]  (.A(addr_0[7]), .B(addr_c6), .Y(addr_n7));
    AX1 \addr_RNO[6]  (.A(addr_c4), .B(addr_0[5]), .C(addr_0[6]), .Y(
        addr_n6));
    XNOR2 \addr_RNO[3]  (.A(addr_0[3]), .B(addr_c2), .Y(addr_n3));
    XOR2 \addr_RNO[1]  (.A(addr_0[1]), .B(addr_0[0]), .Y(addr_n1));
    VCC VCC_i (.Y(VCC));
    DFN0C0 \addr[3]  (.D(addr_n3), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[3]));
    DFN0C0 \addr[8]  (.D(addr_n8), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[8]));
    INV \addr_RNO[0]  (.A(addr_0[0]), .Y(\un1_noise_addr_0_i[0] ));
    OR3B \addr_RNI5BI51[4]  (.A(addr_0[3]), .B(addr_0[4]), .C(addr_c2), 
        .Y(addr_c4));
    DFN0C0 \addr[9]  (.D(addr_n9), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[9]));
    XOR2 \addr_RNO[9]  (.A(addr_0[9]), .B(addr_c8), .Y(addr_n9));
    OR3C \addr_RNI0DHM[2]  (.A(addr_0[0]), .B(addr_0[1]), .C(addr_0[2])
        , .Y(addr_c2));
    DFN0C0 \addr[0]  (.D(\un1_noise_addr_0_i[0] ), .CLK(
        s_clk_div4_0_clkout), .CLR(n_acq_change_0_n_rst_n_0), .Q(
        addr_0[0]));
    DFN0C0 \addr[4]  (.D(addr_n4), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[4]));
    DFN0C0 \addr[5]  (.D(addr_n5), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[5]));
    GND GND_i (.Y(GND));
    AX1C \addr_RNO[2]  (.A(addr_0[0]), .B(addr_0[1]), .C(addr_0[2]), 
        .Y(addr_n2));
    AX1C \addr_RNO[11]  (.A(addr_c9), .B(addr_0[10]), .C(addr_0[11]), 
        .Y(addr_n11));
    DFN0C0 \addr[2]  (.D(addr_n2), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[2]));
    XOR2 \addr_RNO[10]  (.A(addr_0[10]), .B(addr_c9), .Y(addr_n10));
    XNOR2 \addr_RNO[5]  (.A(addr_0[5]), .B(addr_c4), .Y(addr_n5));
    OR3B \addr_RNIE9JK1[6]  (.A(addr_0[5]), .B(addr_0[6]), .C(addr_c4), 
        .Y(addr_c6));
    DFN0C0 \addr[10]  (.D(addr_n10), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n_0), .Q(addr_0[10]));
    DFN0C0 \addr[7]  (.D(addr_n7), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[7]));
    AX1 \addr_RNO[4]  (.A(addr_c2), .B(addr_0[3]), .C(addr_0[4]), .Y(
        addr_n4));
    NOR3B \addr_RNIR7K32[8]  (.A(addr_0[7]), .B(addr_0[8]), .C(addr_c6)
        , .Y(addr_c8));
    DFN0C0 \addr[1]  (.D(addr_n1), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .Q(addr_0[1]));
    AX1 \addr_RNO[8]  (.A(addr_c6), .B(addr_0[7]), .C(addr_0[8]), .Y(
        addr_n8));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR2B \addr_RNI3N4B2[9]  (.A(addr_0[9]), .B(addr_c8), .Y(addr_c9));
    
endmodule


module noiseclk(
       n_divnum,
       top_code_0_n_load,
       GLA,
       s_clk_div4_0_clkout,
       noiseclkctrl_0_en,
       n_acq_change_0_n_acq_start,
       n_acq_change_0_n_rst_n_0
    );
input  [9:0] n_divnum;
input  top_code_0_n_load;
input  GLA;
output s_clk_div4_0_clkout;
input  noiseclkctrl_0_en;
input  n_acq_change_0_n_acq_start;
input  n_acq_change_0_n_rst_n_0;

    wire N_12, \count[1]_net_1 , \count[0]_net_1 , N_4, 
        \count[3]_net_1 , \DWACT_FINC_E[0] , count_0_sqmuxa_1_0_net_1, 
        en_net_1, ADD_5x5_medium_area_I8_Y_0, N87, 
        ADD_5x5_medium_area_I8_un1_Y_0, N88, clkout8_NE_2, clkout8_3_i, 
        clkout8_4_i, clkout8_1_i, clkout8_NE_1, \count[2]_net_1 , 
        \datahalf[2]_net_1 , clkout8_0_i, N96, N94, clkout_1_sqmuxa, 
        I_11, clkout8_NE_i, \dataall_1[4] , N_43, clkout_6, N83, 
        ADD_5x5_medium_area_I9_un1_Y, \dataall_1[0] , \dataall_1[1] , 
        \dataall_1[2] , \dataall_1[3] , \datahalf[0]_net_1 , 
        \datahalf[1]_net_1 , \datahalf[3]_net_1 , \datahalf[4]_net_1 , 
        \count[4]_net_1 , clkout9, \count_6[1] , I_5_2, \count_6[2] , 
        I_9_2, \count_6[3] , I_13_2, \count_6[4] , I_20_2, 
        \count_6[0] , clkout_RNO_net_1, \dataall[0]_net_1 , 
        \dataall[1]_net_1 , \dataall[2]_net_1 , \dataall[3]_net_1 , 
        \dataall[4]_net_1 , N_9, N_13, N_12_0, N_11, N_8, N_10, N_9_0, 
        N_7, N_4_0, N_5, N_6, GND, VCC, GND_0, VCC_0;
    
    AX1D dataall_1_ADD_5x5_medium_area_I12_Y_0 (.A(
        ADD_5x5_medium_area_I9_un1_Y), .B(N87), .C(N88), .Y(
        \dataall_1[3] ));
    XOR3 dataall_1_ADD_5x5_medium_area_I11_Y_0 (.A(n_divnum[2]), .B(
        n_divnum[7]), .C(N94), .Y(\dataall_1[2] ));
    OA1A un1_count_0_I_6 (.A(\count[3]_net_1 ), .B(\dataall[3]_net_1 ), 
        .C(N_5), .Y(N_9_0));
    AO1C un1_count_0_I_7 (.A(\count[2]_net_1 ), .B(\dataall[2]_net_1 ), 
        .C(N_4_0), .Y(N_10));
    NOR2B \datahalf_RNIMOT42[2]  (.A(clkout8_NE_2), .B(clkout8_NE_1), 
        .Y(clkout8_NE_i));
    NOR2B dataall_1_ADD_5x5_medium_area_I2_CO1 (.A(n_divnum[7]), .B(
        n_divnum[2]), .Y(N87));
    DFN1E1 \dataall[4]  (.D(\dataall_1[4] ), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\dataall[4]_net_1 ));
    DFN1 \count[1]  (.D(\count_6[1] ), .CLK(GLA), .Q(\count[1]_net_1 ));
    DFN1E1 \datahalf[1]  (.D(n_divnum[1]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\datahalf[1]_net_1 ));
    DFN1 \count[0]  (.D(\count_6[0] ), .CLK(GLA), .Q(\count[0]_net_1 ));
    AND3 un3_count_I_16 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(\DWACT_FINC_E[0] ));
    MX2 clkout_RNO_0 (.A(clkout_6), .B(s_clk_div4_0_clkout), .S(
        clkout_1_sqmuxa), .Y(N_43));
    NOR3A clkout_RNO_2 (.A(I_11), .B(clkout8_NE_i), .C(en_net_1), .Y(
        clkout_1_sqmuxa));
    XOR3 dataall_1_ADD_5x5_medium_area_I13_Y_0 (.A(n_divnum[4]), .B(
        n_divnum[9]), .C(N96), .Y(\dataall_1[4] ));
    OR2A un1_count_0_I_1 (.A(\dataall[1]_net_1 ), .B(\count[1]_net_1 ), 
        .Y(N_4_0));
    XNOR2 \datahalf_RNI09PD[3]  (.A(\datahalf[3]_net_1 ), .B(
        \count[3]_net_1 ), .Y(clkout8_3_i));
    XA1 dataall_1_ADD_5x5_medium_area_I8_un1_Y_0 (.A(n_divnum[2]), .B(
        n_divnum[7]), .C(N88), .Y(ADD_5x5_medium_area_I8_un1_Y_0));
    NOR3A \count_RNO[2]  (.A(I_9_2), .B(clkout9), .C(
        count_0_sqmuxa_1_0_net_1), .Y(\count_6[2] ));
    VCC VCC_i (.Y(VCC));
    NOR3A \count_RNO[4]  (.A(I_20_2), .B(clkout9), .C(
        count_0_sqmuxa_1_0_net_1), .Y(\count_6[4] ));
    NOR2B clkout_RNO (.A(n_acq_change_0_n_rst_n_0), .B(N_43), .Y(
        clkout_RNO_net_1));
    OR2A count_0_sqmuxa_1_0 (.A(n_acq_change_0_n_rst_n_0), .B(en_net_1)
        , .Y(count_0_sqmuxa_1_0_net_1));
    NOR2 \datahalf_RNIOJE25[2]  (.A(I_11), .B(clkout8_NE_i), .Y(
        clkout9));
    OA1A un1_count_0_I_10 (.A(N_8), .B(N_10), .C(N_9_0), .Y(N_13));
    NOR3C \datahalf_RNIUMB91[1]  (.A(clkout8_3_i), .B(clkout8_4_i), .C(
        clkout8_1_i), .Y(clkout8_NE_2));
    XOR2 un3_count_I_5 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), .Y(
        I_5_2));
    DFN1E1 \dataall[0]  (.D(\dataall_1[0] ), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\dataall[0]_net_1 ));
    NOR2A un1_count_0_I_3 (.A(\dataall[0]_net_1 ), .B(\count[0]_net_1 )
        , .Y(N_6));
    NOR3A \count_RNO[3]  (.A(I_13_2), .B(clkout9), .C(
        count_0_sqmuxa_1_0_net_1), .Y(\count_6[3] ));
    DFN1E1 \dataall[2]  (.D(\dataall_1[2] ), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\dataall[2]_net_1 ));
    NOR2B dataall_1_ADD_5x5_medium_area_I0_CO1 (.A(n_divnum[5]), .B(
        n_divnum[0]), .Y(N83));
    AO1B dataall_1_ADD_5x5_medium_area_I8_Y (.A(
        ADD_5x5_medium_area_I8_un1_Y_0), .B(N94), .C(
        ADD_5x5_medium_area_I8_Y_0), .Y(N96));
    XA1 dataall_1_ADD_5x5_medium_area_I9_un1_Y (.A(n_divnum[2]), .B(
        n_divnum[7]), .C(N94), .Y(ADD_5x5_medium_area_I9_un1_Y));
    NOR3A \count_RNO[1]  (.A(I_5_2), .B(clkout9), .C(
        count_0_sqmuxa_1_0_net_1), .Y(\count_6[1] ));
    XOR2 un3_count_I_9 (.A(N_12), .B(\count[2]_net_1 ), .Y(I_9_2));
    XNOR2 \datahalf_RNIQSOD[0]  (.A(\datahalf[0]_net_1 ), .B(
        \count[0]_net_1 ), .Y(clkout8_0_i));
    DFN1 \count[2]  (.D(\count_6[2] ), .CLK(GLA), .Q(\count[2]_net_1 ));
    OR2B en (.A(n_acq_change_0_n_acq_start), .B(noiseclkctrl_0_en), .Y(
        en_net_1));
    OR2A un1_count_0_I_8 (.A(\count[4]_net_1 ), .B(\dataall[4]_net_1 ), 
        .Y(N_11));
    AO1C un1_count_0_I_5 (.A(\dataall[1]_net_1 ), .B(\count[1]_net_1 ), 
        .C(N_6), .Y(N_8));
    OR2A un1_count_0_I_2 (.A(\count[2]_net_1 ), .B(\dataall[2]_net_1 ), 
        .Y(N_5));
    DFN1 clkout (.D(clkout_RNO_net_1), .CLK(GLA), .Q(
        s_clk_div4_0_clkout));
    AO1C un1_count_0_I_9 (.A(\count[3]_net_1 ), .B(\dataall[3]_net_1 ), 
        .C(N_7), .Y(N_12_0));
    GND GND_i (.Y(GND));
    NOR2B un3_count_I_19 (.A(\count[3]_net_1 ), .B(\DWACT_FINC_E[0] ), 
        .Y(N_4));
    AND3 un3_count_I_12 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(N_9));
    DFN1E1 \dataall[1]  (.D(\dataall_1[1] ), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\dataall[1]_net_1 ));
    OR3A \count_RNO[0]  (.A(\count[0]_net_1 ), .B(clkout9), .C(
        count_0_sqmuxa_1_0_net_1), .Y(\count_6[0] ));
    NOR2B un3_count_I_8 (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .Y(N_12));
    DFN1E1 \datahalf[0]  (.D(n_divnum[0]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\datahalf[0]_net_1 ));
    OR2A un1_count_0_I_4 (.A(\dataall[4]_net_1 ), .B(\count[4]_net_1 ), 
        .Y(N_7));
    XA1A \datahalf_RNIO1IR[2]  (.A(\count[2]_net_1 ), .B(
        \datahalf[2]_net_1 ), .C(clkout8_0_i), .Y(clkout8_NE_1));
    NOR2 clkout_RNO_1 (.A(s_clk_div4_0_clkout), .B(en_net_1), .Y(
        clkout_6));
    XOR3 dataall_1_ADD_5x5_medium_area_I10_Y_0 (.A(n_divnum[1]), .B(
        n_divnum[6]), .C(N83), .Y(\dataall_1[1] ));
    DFN1 \count[3]  (.D(\count_6[3] ), .CLK(GLA), .Q(\count[3]_net_1 ));
    DFN1E1 \datahalf[4]  (.D(n_divnum[4]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\datahalf[4]_net_1 ));
    XNOR2 \datahalf_RNI2DPD[4]  (.A(\datahalf[4]_net_1 ), .B(
        \count[4]_net_1 ), .Y(clkout8_4_i));
    XOR2 dataall_1_ADD_5x5_medium_area_I3_S_0 (.A(n_divnum[8]), .B(
        n_divnum[3]), .Y(N88));
    XOR2 un3_count_I_20 (.A(N_4), .B(\count[4]_net_1 ), .Y(I_20_2));
    OA1 un1_count_0_I_11 (.A(N_13), .B(N_12_0), .C(N_11), .Y(I_11));
    XNOR2 \datahalf_RNIS0PD[1]  (.A(\datahalf[1]_net_1 ), .B(
        \count[1]_net_1 ), .Y(clkout8_1_i));
    MIN3 dataall_1_ADD_5x5_medium_area_I8_Y_0 (.A(n_divnum[3]), .B(
        n_divnum[8]), .C(N87), .Y(ADD_5x5_medium_area_I8_Y_0));
    XOR2 dataall_1_ADD_5x5_medium_area_I0_S_0 (.A(n_divnum[5]), .B(
        n_divnum[0]), .Y(\dataall_1[0] ));
    DFN1E1 \datahalf[2]  (.D(n_divnum[2]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\datahalf[2]_net_1 ));
    DFN1E1 \dataall[3]  (.D(\dataall_1[3] ), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\dataall[3]_net_1 ));
    MAJ3 dataall_1_ADD_5x5_medium_area_I7_Y (.A(n_divnum[1]), .B(
        n_divnum[6]), .C(N83), .Y(N94));
    DFN1 \count[4]  (.D(\count_6[4] ), .CLK(GLA), .Q(\count[4]_net_1 ));
    XOR2 un3_count_I_13 (.A(N_9), .B(\count[3]_net_1 ), .Y(I_13_2));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    DFN1E1 \datahalf[3]  (.D(n_divnum[3]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\datahalf[3]_net_1 ));
    
endmodule


module noiseclkctrl(
       n_acqnum,
       top_code_0_n_load,
       GLA,
       n_acq_change_0_n_rst_n,
       s_clk_div4_0_clkout,
       noiseclkctrl_0_en
    );
input  [11:0] n_acqnum;
input  top_code_0_n_load;
input  GLA;
input  n_acq_change_0_n_rst_n;
input  s_clk_div4_0_clkout;
output noiseclkctrl_0_en;

    wire count_c2, \count[0]_net_1 , \count[1]_net_1 , 
        \count[2]_net_1 , count_c4, \count[3]_net_1 , \count[4]_net_1 , 
        count_c6, \count[5]_net_1 , \count[6]_net_1 , count_c8, 
        \count[7]_net_1 , \count[8]_net_1 , count_c9, \count[9]_net_1 , 
        en_RNO_0, counte, count_n1, \count_RNO_1[0] , count_n2, 
        count_n3, count_n4, count_n5, count_n6, count_n7, count_n8, 
        count_n9, count_n10, \count[10]_net_1 , count_n11, 
        \count[11]_net_1 , \data[0]_net_1 , \data[1]_net_1 , 
        \data[2]_net_1 , \data[3]_net_1 , \data[4]_net_1 , 
        \data[5]_net_1 , \data[6]_net_1 , \data[7]_net_1 , 
        \data[8]_net_1 , \data[9]_net_1 , \data[10]_net_1 , 
        \data[11]_net_1 , \DWACT_COMP0_E[1] , \DWACT_COMP0_E[2] , 
        \DWACT_COMP0_E[0] , \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] , 
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] , \ACT_LT4_E[3] , 
        \ACT_LT4_E[6] , \ACT_LT4_E[10] , \ACT_LT4_E[7] , 
        \ACT_LT4_E[8] , \ACT_LT4_E[5] , \ACT_LT4_E[4] , \ACT_LT4_E[0] , 
        \ACT_LT4_E[1] , \ACT_LT4_E[2] , \ACT_LT3_E[3] , \ACT_LT3_E[4] , 
        \ACT_LT3_E[5] , \ACT_LT3_E[0] , \ACT_LT3_E[1] , \ACT_LT3_E[2] , 
        \DWACT_BL_EQUAL_0_E[2] , \DWACT_BL_EQUAL_0_E[1] , 
        \DWACT_BL_EQUAL_0_E[0] , N_37, N_36, N_35, N_32, N_34, N_33, 
        N_31, N_28, N_29, N_30, \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] , 
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] , \DWACT_BL_EQUAL_0_E[4] , 
        \DWACT_BL_EQUAL_0_E[3] , \DWACT_BL_EQUAL_0_E_0[0] , 
        \DWACT_BL_EQUAL_0_E_0[1] , \DWACT_BL_EQUAL_0_E_0[2] , GND, VCC, 
        GND_0, VCC_0;
    
    NOR2A un1_count_0_I_62 (.A(\count[2]_net_1 ), .B(\data[2]_net_1 ), 
        .Y(\ACT_LT4_E[7] ));
    AND2A un1_count_0_I_57 (.A(\data[1]_net_1 ), .B(\count[1]_net_1 ), 
        .Y(\ACT_LT4_E[2] ));
    AO1 un1_count_0_I_72 (.A(\DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ), .B(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ), .C(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ), .Y(\DWACT_COMP0_E[2] ));
    AND3 un1_count_0_I_6 (.A(\DWACT_BL_EQUAL_0_E_0[0] ), .B(
        \DWACT_BL_EQUAL_0_E_0[1] ), .C(\DWACT_BL_EQUAL_0_E_0[2] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ));
    OA1 un1_count_0_I_27 (.A(N_37), .B(N_36), .C(N_35), .Y(
        \DWACT_COMP0_E[0] ));
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[5]_net_1 ));
    AND2 un1_count_0_I_7 (.A(\DWACT_BL_EQUAL_0_E[4] ), .B(
        \DWACT_BL_EQUAL_0_E[3] ), .Y(
        \DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ));
    OR2A un1_count_0_I_59 (.A(\data[2]_net_1 ), .B(\count[2]_net_1 ), 
        .Y(\ACT_LT4_E[4] ));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[1]_net_1 ));
    DFN1E1 \data[3]  (.D(n_acqnum[3]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[3]_net_1 ));
    NOR2B \count_RNI5GE52[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_c9));
    DFN1E1C0 \count[10]  (.D(count_n10), .CLK(s_clk_div4_0_clkout), 
        .CLR(n_acq_change_0_n_rst_n), .E(counte), .Q(\count[10]_net_1 )
        );
    DFN1P0 \count[0]  (.D(\count_RNO_1[0] ), .CLK(s_clk_div4_0_clkout), 
        .PRE(n_acq_change_0_n_rst_n), .Q(\count[0]_net_1 ));
    DFN1E1 \data[5]  (.D(n_acqnum[5]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[5]_net_1 ));
    OR2A un1_count_0_I_63 (.A(\count[3]_net_1 ), .B(\data[3]_net_1 ), 
        .Y(\ACT_LT4_E[8] ));
    AO1C un1_count_0_I_21 (.A(\data[8]_net_1 ), .B(\count[8]_net_1 ), 
        .C(N_30), .Y(N_32));
    AND2A un1_count_0_I_47 (.A(\data[6]_net_1 ), .B(\count[6]_net_1 ), 
        .Y(\ACT_LT3_E[5] ));
    XOR2 \count_RNO[7]  (.A(count_c6), .B(\count[7]_net_1 ), .Y(
        count_n7));
    NOR2A un1_count_0_I_60 (.A(\data[3]_net_1 ), .B(\count[3]_net_1 ), 
        .Y(\ACT_LT4_E[5] ));
    XNOR2 un1_count_0_I_1 (.A(\count[11]_net_1 ), .B(\data[11]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E[4] ));
    AX1C \count_RNO[2]  (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(count_n2));
    DFN1E1 \data[9]  (.D(n_acqnum[9]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[9]_net_1 ));
    XOR2 \count_RNO[9]  (.A(count_c8), .B(\count[9]_net_1 ), .Y(
        count_n9));
    DFN1E1 \data[2]  (.D(n_acqnum[2]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[2]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1 \data[6]  (.D(n_acqnum[6]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[6]_net_1 ));
    AX1C \count_RNO[4]  (.A(\count[3]_net_1 ), .B(count_c2), .C(
        \count[4]_net_1 ), .Y(count_n4));
    DFN1E1C0 \count[8]  (.D(count_n8), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[8]_net_1 ));
    DFN1E1 \data[7]  (.D(n_acqnum[7]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[7]_net_1 ));
    DFN1E1 \data[10]  (.D(n_acqnum[10]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\data[10]_net_1 ));
    XNOR2 un1_count_0_I_36 (.A(\count[6]_net_1 ), .B(\data[6]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E[2] ));
    NOR2B en_RNO (.A(noiseclkctrl_0_en), .B(counte), .Y(en_RNO_0));
    AOI1A un1_count_0_I_64 (.A(\ACT_LT4_E[7] ), .B(\ACT_LT4_E[8] ), .C(
        \ACT_LT4_E[5] ), .Y(\ACT_LT4_E[10] ));
    XOR2 \count_RNO[10]  (.A(count_c9), .B(\count[10]_net_1 ), .Y(
        count_n10));
    AOI1A un1_count_0_I_65 (.A(\ACT_LT4_E[3] ), .B(\ACT_LT4_E[6] ), .C(
        \ACT_LT4_E[10] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[2] ));
    DFN1E1 \data[0]  (.D(n_acqnum[0]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[0]_net_1 ));
    NOR3C \count_RNINDPK[2]  (.A(\count[0]_net_1 ), .B(
        \count[1]_net_1 ), .C(\count[2]_net_1 ), .Y(count_c2));
    DFN1E1 \data[11]  (.D(n_acqnum[11]), .CLK(GLA), .E(
        top_code_0_n_load), .Q(\data[11]_net_1 ));
    XNOR2 un1_count_0_I_3 (.A(\count[9]_net_1 ), .B(\data[9]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E_0[2] ));
    XOR2 \count_RNO[3]  (.A(count_c2), .B(\count[3]_net_1 ), .Y(
        count_n3));
    DFN1E1C0 \count[11]  (.D(count_n11), .CLK(s_clk_div4_0_clkout), 
        .CLR(n_acq_change_0_n_rst_n), .E(counte), .Q(\count[11]_net_1 )
        );
    DFN1E1 \data[8]  (.D(n_acqnum[8]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[8]_net_1 ));
    AX1C \count_RNO[8]  (.A(\count[7]_net_1 ), .B(count_c6), .C(
        \count[8]_net_1 ), .Y(count_n8));
    XOR2 \count_RNO[5]  (.A(count_c4), .B(\count[5]_net_1 ), .Y(
        count_n5));
    XOR2 \count_RNO[1]  (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .Y(count_n1));
    AX1C \count_RNO[11]  (.A(\count[10]_net_1 ), .B(count_c9), .C(
        \count[11]_net_1 ), .Y(count_n11));
    OR2A un1_count_0_I_56 (.A(\data[1]_net_1 ), .B(\count[1]_net_1 ), 
        .Y(\ACT_LT4_E[1] ));
    OA1A un1_count_0_I_26 (.A(N_32), .B(N_34), .C(N_33), .Y(N_37));
    DFN1E1 \data[4]  (.D(n_acqnum[4]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[4]_net_1 ));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[2]_net_1 ));
    DFN1P0 en (.D(en_RNO_0), .CLK(s_clk_div4_0_clkout), .PRE(
        n_acq_change_0_n_rst_n), .Q(noiseclkctrl_0_en));
    AND2 un1_count_0_I_8 (.A(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[1] ), 
        .B(\DWACT_BL_EQUAL_0_DWACT_ANDTREE_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    XNOR2 un1_count_0_I_5 (.A(\count[8]_net_1 ), .B(\data[8]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E_0[1] ));
    OA1A un1_count_0_I_22 (.A(\count[10]_net_1 ), .B(\data[10]_net_1 ), 
        .C(N_29), .Y(N_33));
    XNOR2 un1_count_0_I_2 (.A(\count[7]_net_1 ), .B(\data[7]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E_0[0] ));
    NOR3C \count_RNIPDIG1[6]  (.A(\count[5]_net_1 ), .B(count_c4), .C(
        \count[6]_net_1 ), .Y(count_c6));
    OR2A un1_count_0_I_18 (.A(\count[9]_net_1 ), .B(\data[9]_net_1 ), 
        .Y(N_29));
    GND GND_i (.Y(GND));
    DFN1E1C0 \count[9]  (.D(count_n9), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[9]_net_1 ));
    AO1 un1_count_0_I_77 (.A(\DWACT_COMP0_E[1] ), .B(
        \DWACT_COMP0_E[2] ), .C(\DWACT_COMP0_E[0] ), .Y(counte));
    AX1C \count_RNO[6]  (.A(\count[5]_net_1 ), .B(count_c4), .C(
        \count[6]_net_1 ), .Y(count_n6));
    XOR2 \count_RNO[0]  (.A(counte), .B(\count[0]_net_1 ), .Y(
        \count_RNO_1[0] ));
    OR2A un1_count_0_I_46 (.A(\data[6]_net_1 ), .B(\count[6]_net_1 ), 
        .Y(\ACT_LT3_E[4] ));
    AO1C un1_count_0_I_23 (.A(\count[9]_net_1 ), .B(\data[9]_net_1 ), 
        .C(N_28), .Y(N_34));
    NOR2A un1_count_0_I_42 (.A(\data[4]_net_1 ), .B(\count[4]_net_1 ), 
        .Y(\ACT_LT3_E[0] ));
    NOR2A un1_count_0_I_61 (.A(\ACT_LT4_E[4] ), .B(\ACT_LT4_E[5] ), .Y(
        \ACT_LT4_E[6] ));
    XNOR2 un1_count_0_I_4 (.A(\count[10]_net_1 ), .B(\data[10]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E[3] ));
    XNOR2 un1_count_0_I_34 (.A(\count[4]_net_1 ), .B(\data[4]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E[0] ));
    XNOR2 un1_count_0_I_35 (.A(\count[5]_net_1 ), .B(\data[5]_net_1 ), 
        .Y(\DWACT_BL_EQUAL_0_E[1] ));
    OR2A un1_count_0_I_20 (.A(\data[11]_net_1 ), .B(\count[11]_net_1 ), 
        .Y(N_31));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[6]_net_1 ));
    OR2A un1_count_0_I_43 (.A(\data[5]_net_1 ), .B(\count[5]_net_1 ), 
        .Y(\ACT_LT3_E[1] ));
    OR2A un1_count_0_I_17 (.A(\data[8]_net_1 ), .B(\count[8]_net_1 ), 
        .Y(N_28));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[3]_net_1 ));
    NOR2A un1_count_0_I_19 (.A(\data[7]_net_1 ), .B(\count[7]_net_1 ), 
        .Y(N_30));
    DFN1E1 \data[1]  (.D(n_acqnum[1]), .CLK(GLA), .E(top_code_0_n_load)
        , .Q(\data[1]_net_1 ));
    NOR2A un1_count_0_I_55 (.A(\data[0]_net_1 ), .B(\count[0]_net_1 ), 
        .Y(\ACT_LT4_E[0] ));
    OR2A un1_count_0_I_24 (.A(\count[11]_net_1 ), .B(\data[11]_net_1 ), 
        .Y(N_35));
    AO1C un1_count_0_I_25 (.A(\count[10]_net_1 ), .B(\data[10]_net_1 ), 
        .C(N_31), .Y(N_36));
    NOR3C \count_RNIMLL21[4]  (.A(\count[3]_net_1 ), .B(count_c2), .C(
        \count[4]_net_1 ), .Y(count_c4));
    AND3 un1_count_0_I_37 (.A(\DWACT_BL_EQUAL_0_E[2] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E[0] ), .Y(
        \DWACT_CMPLE_PO2_DWACT_COMP0_E[1] ));
    AOI1A un1_count_0_I_58 (.A(\ACT_LT4_E[0] ), .B(\ACT_LT4_E[1] ), .C(
        \ACT_LT4_E[2] ), .Y(\ACT_LT4_E[3] ));
    AND2A un1_count_0_I_44 (.A(\data[5]_net_1 ), .B(\count[5]_net_1 ), 
        .Y(\ACT_LT3_E[2] ));
    AOI1A un1_count_0_I_45 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), .C(
        \ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    NOR3C \count_RNI0MFU1[7]  (.A(\count[7]_net_1 ), .B(count_c6), .C(
        \count[8]_net_1 ), .Y(count_c8));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[4]_net_1 ));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(s_clk_div4_0_clkout), .CLR(
        n_acq_change_0_n_rst_n), .E(counte), .Q(\count[7]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    AOI1A un1_count_0_I_48 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), .C(
        \ACT_LT3_E[5] ), .Y(\DWACT_CMPLE_PO2_DWACT_COMP0_E[0] ));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module RAM(
       un1_n_s_change_0,
       addr_0,
       addr,
       MX2_RD_8_inst,
       MX2_RD_10_inst,
       MX2_RD_3_inst,
       MX2_RD_9_inst,
       MX2_RD_1_inst,
       top_code_0_n_rd_en,
       MX2_RD_11_inst,
       MX2_RD_6_inst,
       MX2_RD_7_inst,
       n_acq_change_0_n_acq_start,
       MX2_RD_5_inst,
       MX2_RD_4_inst,
       s_clk_div4_0_clkout,
       RAM_VCC,
       n_acq_change_0_n_rst_n_0,
       n_rdclk,
       RAM_GND,
       MX2_RD_2_inst,
       MX2_RD_0_inst
    );
input  [11:0] un1_n_s_change_0;
input  [11:0] addr_0;
input  [11:0] addr;
output MX2_RD_8_inst;
output MX2_RD_10_inst;
output MX2_RD_3_inst;
output MX2_RD_9_inst;
output MX2_RD_1_inst;
input  top_code_0_n_rd_en;
output MX2_RD_11_inst;
output MX2_RD_6_inst;
output MX2_RD_7_inst;
input  n_acq_change_0_n_acq_start;
output MX2_RD_5_inst;
output MX2_RD_4_inst;
input  s_clk_div4_0_clkout;
input  RAM_VCC;
input  n_acq_change_0_n_rst_n_0;
input  n_rdclk;
input  RAM_GND;
output MX2_RD_2_inst;
output MX2_RD_0_inst;

    wire MX2_149_Y, MX2_75_Y, MX2_127_Y, BUFF_16_Y, MX2_140_Y, 
        MX2_14_Y, MX2_147_Y, BUFF_17_Y, MX2_144_Y, QX_TEMPR10_5_net, 
        QX_TEMPR11_5_net, BUFF_12_Y, BLKB_EN_2_net, ENABLE_ADDRB_2_net, 
        WEBP, MX2_13_Y, QX_TEMPR8_8_net, QX_TEMPR9_8_net, BUFF_1_Y, 
        BLKB_EN_5_net, ENABLE_ADDRB_5_net, MX2_1_Y, QX_TEMPR10_6_net, 
        QX_TEMPR11_6_net, MX2_162_Y, MX2_22_Y, MX2_111_Y, BUFF_18_Y, 
        ADDRB_FF2_0_net, MX2_126_Y, QX_TEMPR6_10_net, QX_TEMPR7_10_net, 
        BUFF_6_Y, BLKB_EN_10_net, ENABLE_ADDRB_10_net, ADDRB_FF2_1_net, 
        MX2_85_Y, QX_TEMPR14_3_net, QX_TEMPR15_3_net, BUFF_13_Y, 
        BLKA_EN_8_net, ENABLE_ADDRA_8_net, WEAP, MX2_16_Y, MX2_3_Y, 
        MX2_167_Y, BUFF_5_Y, MX2_165_Y, MX2_34_Y, BUFF_0_Y, MX2_122_Y, 
        MX2_118_Y, MX2_94_Y, MX2_129_Y, MX2_17_Y, BUFF_3_Y, 
        ENABLE_ADDRA_12_net, NOR2_2_Y, AND2_1_Y, BLKA_EN_13_net, 
        ENABLE_ADDRA_13_net, MX2_137_Y, QX_TEMPR8_4_net, 
        QX_TEMPR9_4_net, BUFF_14_Y, BUFF_11_Y, QX_TEMPR7_0_net, 
        QX_TEMPR7_1_net, QX_TEMPR7_2_net, QX_TEMPR7_3_net, 
        QX_TEMPR7_4_net, QX_TEMPR7_5_net, QX_TEMPR7_6_net, 
        QX_TEMPR7_7_net, QX_TEMPR7_8_net, QX_TEMPR7_9_net, 
        QX_TEMPR7_11_net, RAM_R7C0_RD12, RAM_R7C0_RD13, RAM_R7C0_RD14, 
        RAM_R7C0_RD15, RAM_R7C0_RD16, RAM_R7C0_RD17, BLKB_EN_7_net, 
        BLKA_EN_7_net, MX2_18_Y, QX_TEMPR12_10_net, QX_TEMPR13_10_net, 
        BUFF_7_Y, MX2_138_Y, MX2_19_Y, MX2_99_Y, BLKB_EN_3_net, 
        ENABLE_ADDRB_3_net, MX2_161_Y, MX2_108_Y, BUFF_15_Y, 
        ENABLE_ADDRA_5_net, AND2A_2_Y, AND2A_0_Y, MX2_47_Y, 
        QX_TEMPR10_10_net, QX_TEMPR11_10_net, QX_TEMPR6_3_net, 
        BLKA_EN_6_net, ENABLE_ADDRA_6_net, AND2_0_Y, NOR2_3_Y, 
        ENABLE_ADDRA_3_net, AND2_2_Y, NOR2_1_Y, MX2_73_Y, MX2_21_Y, 
        MX2_101_Y, QX_TEMPR8_7_net, QX_TEMPR9_7_net, BUFF_4_Y, 
        MX2_81_Y, MX2_135_Y, MX2_28_Y, BUFF_10_Y, MX2_89_Y, MX2_87_Y, 
        QX_TEMPR2_10_net, QX_TEMPR3_10_net, MX2_74_Y, QX_TEMPR14_9_net, 
        QX_TEMPR15_9_net, MX2_39_Y, MX2_53_Y, MX2_8_Y, MX2_12_Y, 
        QX_TEMPR8_5_net, QX_TEMPR9_5_net, MX2_64_Y, QX_TEMPR0_0_net, 
        QX_TEMPR1_0_net, ENABLE_ADDRB_8_net, NOR2_0_Y, AND2A_5_Y, 
        MX2_103_Y, MX2_59_Y, MX2_120_Y, MX2_145_Y, MX2_4_Y, MX2_104_Y, 
        QX_TEMPR10_0_net, QX_TEMPR10_1_net, QX_TEMPR10_2_net, 
        QX_TEMPR10_3_net, QX_TEMPR10_4_net, QX_TEMPR10_7_net, 
        QX_TEMPR10_8_net, QX_TEMPR10_9_net, QX_TEMPR10_11_net, 
        RAM_R10C0_RD12, RAM_R10C0_RD13, RAM_R10C0_RD14, RAM_R10C0_RD15, 
        RAM_R10C0_RD16, RAM_R10C0_RD17, BLKA_EN_10_net, MX2_50_Y, 
        MX2_97_Y, MX2_43_Y, QX_TEMPR11_2_net, BUFF_2_Y, MX2_79_Y, 
        QX_TEMPR14_11_net, QX_TEMPR15_11_net, QX_TEMPR3_0_net, 
        QX_TEMPR3_1_net, QX_TEMPR3_2_net, QX_TEMPR3_3_net, 
        QX_TEMPR3_4_net, QX_TEMPR3_5_net, QX_TEMPR3_6_net, 
        QX_TEMPR3_7_net, QX_TEMPR3_8_net, QX_TEMPR3_9_net, 
        QX_TEMPR3_11_net, RAM_R3C0_RD12, RAM_R3C0_RD13, RAM_R3C0_RD14, 
        RAM_R3C0_RD15, RAM_R3C0_RD16, RAM_R3C0_RD17, BLKA_EN_3_net, 
        QX_TEMPR0_9_net, QX_TEMPR1_9_net, BLKB_EN_1_net, 
        ENABLE_ADDRB_1_net, ENABLE_ADDRA_4_net, ENABLE_ADDRA_9_net, 
        AND2A_1_Y, QX_TEMPR6_0_net, QX_TEMPR6_1_net, QX_TEMPR6_2_net, 
        QX_TEMPR6_4_net, QX_TEMPR6_5_net, QX_TEMPR6_6_net, 
        QX_TEMPR6_7_net, QX_TEMPR6_8_net, QX_TEMPR6_9_net, 
        QX_TEMPR6_11_net, RAM_R6C0_RD12, RAM_R6C0_RD13, RAM_R6C0_RD14, 
        RAM_R6C0_RD15, RAM_R6C0_RD16, RAM_R6C0_RD17, BLKB_EN_6_net, 
        MX2_151_Y, QX_TEMPR2_2_net, MX2_69_Y, QX_TEMPR4_2_net, 
        QX_TEMPR5_2_net, ADDRB_FF2_2_net, MX2_106_Y, QX_TEMPR14_5_net, 
        QX_TEMPR15_5_net, ADDRB_FF2_3_net, MX2_46_Y, MX2_78_Y, 
        MX2_31_Y, QX_TEMPR2_3_net, AND2A_6_Y, BLKA_EN_11_net, 
        ENABLE_ADDRA_11_net, MX2_153_Y, QX_TEMPR4_9_net, 
        QX_TEMPR5_9_net, MX2_55_Y, QX_TEMPR8_2_net, QX_TEMPR9_2_net, 
        QX_TEMPR1_1_net, QX_TEMPR1_2_net, QX_TEMPR1_3_net, 
        QX_TEMPR1_4_net, QX_TEMPR1_5_net, QX_TEMPR1_6_net, 
        QX_TEMPR1_7_net, QX_TEMPR1_8_net, QX_TEMPR1_10_net, 
        QX_TEMPR1_11_net, RAM_R1C0_RD12, RAM_R1C0_RD13, RAM_R1C0_RD14, 
        RAM_R1C0_RD15, RAM_R1C0_RD16, RAM_R1C0_RD17, BLKA_EN_1_net, 
        MX2_128_Y, QX_TEMPR8_10_net, QX_TEMPR9_10_net, 
        ENABLE_ADDRA_2_net, AND2A_4_Y, MX2_48_Y, MX2_113_Y, MX2_136_Y, 
        QX_TEMPR11_9_net, ENABLE_ADDRA_10_net, MX2_24_Y, 
        QX_TEMPR12_6_net, QX_TEMPR13_6_net, AND2A_3_Y, MX2_139_Y, 
        MX2_84_Y, MX2_130_Y, MX2_142_Y, MX2_70_Y, MX2_134_Y, 
        QX_TEMPR14_4_net, QX_TEMPR15_4_net, MX2_156_Y, QX_TEMPR4_8_net, 
        QX_TEMPR5_8_net, MX2_102_Y, MX2_71_Y, BUFF_8_Y, MX2_37_Y, 
        QX_TEMPR2_6_net, MX2_29_Y, QX_TEMPR12_4_net, QX_TEMPR13_4_net, 
        MX2_51_Y, MX2_83_Y, MX2_33_Y, MX2_42_Y, QX_TEMPR0_6_net, 
        ENABLE_ADDRA_14_net, MX2_160_Y, QX_TEMPR12_5_net, 
        QX_TEMPR13_5_net, QX_TEMPR15_0_net, QX_TEMPR15_1_net, 
        QX_TEMPR15_2_net, QX_TEMPR15_6_net, QX_TEMPR15_7_net, 
        QX_TEMPR15_8_net, QX_TEMPR15_10_net, RAM_R15C0_RD12, 
        RAM_R15C0_RD13, RAM_R15C0_RD14, RAM_R15C0_RD15, RAM_R15C0_RD16, 
        RAM_R15C0_RD17, BLKB_EN_15_net, BLKA_EN_15_net, MX2_164_Y, 
        QX_TEMPR12_11_net, QX_TEMPR13_11_net, MX2_10_Y, 
        ENABLE_ADDRB_7_net, MX2_77_Y, MX2_163_Y, MX2_157_Y, 
        ENABLE_ADDRB_0_net, QX_TEMPR11_0_net, QX_TEMPR11_1_net, 
        QX_TEMPR11_3_net, QX_TEMPR11_4_net, QX_TEMPR11_7_net, 
        QX_TEMPR11_8_net, QX_TEMPR11_11_net, RAM_R11C0_RD12, 
        RAM_R11C0_RD13, RAM_R11C0_RD14, RAM_R11C0_RD15, RAM_R11C0_RD16, 
        RAM_R11C0_RD17, BLKB_EN_11_net, MX2_93_Y, QX_TEMPR8_11_net, 
        QX_TEMPR9_11_net, MX2_9_Y, MX2_119_Y, MX2_57_Y, MX2_116_Y, 
        MX2_98_Y, MX2_27_Y, QX_TEMPR13_0_net, QX_TEMPR13_1_net, 
        QX_TEMPR13_2_net, QX_TEMPR13_3_net, QX_TEMPR13_7_net, 
        QX_TEMPR13_8_net, QX_TEMPR13_9_net, RAM_R13C0_RD12, 
        RAM_R13C0_RD13, RAM_R13C0_RD14, RAM_R13C0_RD15, RAM_R13C0_RD16, 
        RAM_R13C0_RD17, BLKB_EN_13_net, MX2_152_Y, MX2_65_Y, MX2_67_Y, 
        QX_TEMPR0_2_net, QX_TEMPR14_7_net, QX_TEMPR0_10_net, MX2_96_Y, 
        QX_TEMPR14_10_net, MX2_15_Y, QX_TEMPR4_6_net, QX_TEMPR5_6_net, 
        MX2_107_Y, MX2_112_Y, BUFF_9_Y, MX2_7_Y, ENABLE_ADDRB_4_net, 
        MX2_132_Y, MX2_82_Y, QX_TEMPR0_1_net, MX2_36_Y, 
        QX_TEMPR2_8_net, MX2_124_Y, ENABLE_ADDRB_11_net, AND2A_7_Y, 
        MX2_63_Y, MX2_150_Y, MX2_95_Y, MX2_6_Y, MX2_146_Y, MX2_100_Y, 
        BLKA_EN_9_net, MX2_76_Y, MX2_60_Y, MX2_38_Y, QX_TEMPR14_8_net, 
        MX2_121_Y, MX2_11_Y, MX2_41_Y, MX2_45_Y, MX2_56_Y, 
        ENABLE_ADDRB_15_net, AND2_3_Y, MX2_66_Y, MX2_131_Y, MX2_72_Y, 
        BLKB_EN_8_net, MX2_148_Y, MX2_158_Y, MX2_80_Y, MX2_166_Y, 
        QX_TEMPR8_0_net, QX_TEMPR8_1_net, QX_TEMPR8_3_net, 
        QX_TEMPR8_6_net, QX_TEMPR8_9_net, RAM_R8C0_RD12, RAM_R8C0_RD13, 
        RAM_R8C0_RD14, RAM_R8C0_RD15, RAM_R8C0_RD16, RAM_R8C0_RD17, 
        MX2_92_Y, MX2_125_Y, MX2_40_Y, MX2_20_Y, MX2_52_Y, 
        QX_TEMPR12_1_net, BLKA_EN_4_net, QX_TEMPR14_0_net, 
        QX_TEMPR14_1_net, QX_TEMPR14_2_net, QX_TEMPR14_6_net, 
        RAM_R14C0_RD12, RAM_R14C0_RD13, RAM_R14C0_RD14, RAM_R14C0_RD15, 
        RAM_R14C0_RD16, RAM_R14C0_RD17, BLKB_EN_14_net, BLKA_EN_14_net, 
        MX2_32_Y, MX2_105_Y, MX2_68_Y, ENABLE_ADDRB_6_net, MX2_117_Y, 
        MX2_23_Y, QX_TEMPR4_10_net, QX_TEMPR5_10_net, MX2_2_Y, 
        ENABLE_ADDRB_13_net, MX2_61_Y, QX_TEMPR9_1_net, MX2_62_Y, 
        QX_TEMPR9_3_net, QX_TEMPR4_4_net, QX_TEMPR5_4_net, MX2_26_Y, 
        MX2_109_Y, MX2_133_Y, QX_TEMPR2_0_net, QX_TEMPR2_1_net, 
        QX_TEMPR2_4_net, QX_TEMPR2_5_net, QX_TEMPR2_7_net, 
        QX_TEMPR2_9_net, QX_TEMPR2_11_net, RAM_R2C0_RD12, 
        RAM_R2C0_RD13, RAM_R2C0_RD14, RAM_R2C0_RD15, RAM_R2C0_RD16, 
        RAM_R2C0_RD17, BLKA_EN_2_net, MX2_141_Y, BLKA_EN_0_net, 
        ENABLE_ADDRA_0_net, MX2_143_Y, MX2_0_Y, QX_TEMPR4_5_net, 
        QX_TEMPR5_5_net, MX2_159_Y, MX2_54_Y, MX2_90_Y, 
        QX_TEMPR12_8_net, QX_TEMPR0_7_net, MX2_154_Y, BLKA_EN_5_net, 
        QX_TEMPR9_9_net, MX2_30_Y, MX2_91_Y, QX_TEMPR0_8_net, 
        QX_TEMPR4_0_net, QX_TEMPR5_0_net, ENABLE_ADDRA_7_net, 
        QX_TEMPR4_11_net, QX_TEMPR5_11_net, MX2_110_Y, QX_TEMPR0_5_net, 
        MX2_114_Y, QX_TEMPR12_7_net, MX2_123_Y, ENABLE_ADDRA_1_net, 
        MX2_35_Y, MX2_49_Y, MX2_86_Y, QX_TEMPR9_0_net, QX_TEMPR9_6_net, 
        RAM_R9C0_RD12, RAM_R9C0_RD13, RAM_R9C0_RD14, RAM_R9C0_RD15, 
        RAM_R9C0_RD16, RAM_R9C0_RD17, BLKB_EN_9_net, QX_TEMPR0_3_net, 
        ENABLE_ADDRA_15_net, BLKB_EN_12_net, ENABLE_ADDRB_12_net, 
        MX2_25_Y, MX2_155_Y, MX2_88_Y, MX2_58_Y, QX_TEMPR4_3_net, 
        QX_TEMPR5_3_net, QX_TEMPR0_4_net, ENABLE_ADDRB_9_net, 
        QX_TEMPR4_7_net, QX_TEMPR5_7_net, MX2_115_Y, 
        ENABLE_ADDRB_14_net, QX_TEMPR12_3_net, BLKB_EN_4_net, 
        QX_TEMPR12_2_net, MX2_5_Y, QX_TEMPR4_1_net, RAM_R4C0_RD12, 
        RAM_R4C0_RD13, RAM_R4C0_RD14, RAM_R4C0_RD15, RAM_R4C0_RD16, 
        RAM_R4C0_RD17, QX_TEMPR12_0_net, QX_TEMPR12_9_net, 
        RAM_R12C0_RD12, RAM_R12C0_RD13, RAM_R12C0_RD14, RAM_R12C0_RD15, 
        RAM_R12C0_RD16, RAM_R12C0_RD17, BLKA_EN_12_net, MX2_44_Y, 
        QX_TEMPR0_11_net, RAM_R0C0_RD12, RAM_R0C0_RD13, RAM_R0C0_RD14, 
        RAM_R0C0_RD15, RAM_R0C0_RD16, RAM_R0C0_RD17, BLKB_EN_0_net, 
        QX_TEMPR5_1_net, RAM_R5C0_RD12, RAM_R5C0_RD13, RAM_R5C0_RD14, 
        RAM_R5C0_RD15, RAM_R5C0_RD16, RAM_R5C0_RD17, GND, VCC, GND_0, 
        VCC_0;
    
    NAND2 NAND2_ENABLE_ADDRB_11_inst (.A(AND2_0_Y), .B(AND2A_5_Y), .Y(
        ENABLE_ADDRB_11_net));
    MX2 MX2_52 (.A(QX_TEMPR2_4_net), .B(QX_TEMPR3_4_net), .S(BUFF_14_Y)
        , .Y(MX2_52_Y));
    MX2 MX2_123 (.A(QX_TEMPR12_9_net), .B(QX_TEMPR13_9_net), .S(
        BUFF_6_Y), .Y(MX2_123_Y));
    AND2 AND2_2 (.A(addr_0[9]), .B(addr_0[8]), .Y(AND2_2_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R5C0.mem") )  RAM_R5C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_5_net), .WEN(BLKA_EN_5_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R5C0_RD17), .RD16(RAM_R5C0_RD16), .RD15(
        RAM_R5C0_RD15), .RD14(RAM_R5C0_RD14), .RD13(RAM_R5C0_RD13), 
        .RD12(RAM_R5C0_RD12), .RD11(QX_TEMPR5_11_net), .RD10(
        QX_TEMPR5_10_net), .RD9(QX_TEMPR5_9_net), .RD8(QX_TEMPR5_8_net)
        , .RD7(QX_TEMPR5_7_net), .RD6(QX_TEMPR5_6_net), .RD5(
        QX_TEMPR5_5_net), .RD4(QX_TEMPR5_4_net), .RD3(QX_TEMPR5_3_net), 
        .RD2(QX_TEMPR5_2_net), .RD1(QX_TEMPR5_1_net), .RD0(
        QX_TEMPR5_0_net));
    NOR2 NOR2_2 (.A(addr_0[9]), .B(addr_0[8]), .Y(NOR2_2_Y));
    MX2 MX2_80 (.A(QX_TEMPR0_11_net), .B(QX_TEMPR1_11_net), .S(
        BUFF_7_Y), .Y(MX2_80_Y));
    OR2 ORA_GATE_10_inst (.A(ENABLE_ADDRA_10_net), .B(WEAP), .Y(
        BLKA_EN_10_net));
    OR2 ORA_GATE_0_inst (.A(ENABLE_ADDRA_0_net), .B(WEAP), .Y(
        BLKA_EN_0_net));
    MX2 MX2_132 (.A(QX_TEMPR12_0_net), .B(QX_TEMPR13_0_net), .S(
        BUFF_11_Y), .Y(MX2_132_Y));
    OR2 ORB_GATE_13_inst (.A(ENABLE_ADDRB_13_net), .B(WEBP), .Y(
        BLKB_EN_13_net));
    BUFF BUFF_10 (.A(ADDRB_FF2_2_net), .Y(BUFF_10_Y));
    MX2 MX2_17 (.A(QX_TEMPR2_1_net), .B(QX_TEMPR3_1_net), .S(BUFF_11_Y)
        , .Y(MX2_17_Y));
    MX2 MX2_121 (.A(QX_TEMPR14_6_net), .B(QX_TEMPR15_6_net), .S(
        BUFF_4_Y), .Y(MX2_121_Y));
    MX2 MX2_166 (.A(QX_TEMPR2_11_net), .B(QX_TEMPR3_11_net), .S(
        BUFF_7_Y), .Y(MX2_166_Y));
    MX2 MX2_58 (.A(MX2_11_Y), .B(MX2_5_Y), .S(BUFF_10_Y), .Y(MX2_58_Y));
    MX2 MX2_49 (.A(QX_TEMPR4_1_net), .B(QX_TEMPR5_1_net), .S(BUFF_11_Y)
        , .Y(MX2_49_Y));
    BUFF BUFF_8 (.A(ADDRB_FF2_1_net), .Y(BUFF_8_Y));
    MX2 MX2_21 (.A(MX2_69_Y), .B(MX2_141_Y), .S(BUFF_3_Y), .Y(MX2_21_Y)
        );
    RAM512X18 #( .MEMORYFILE("RAM_R0C0.mem") )  RAM_R0C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_0_net), .WEN(BLKA_EN_0_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R0C0_RD17), .RD16(RAM_R0C0_RD16), .RD15(
        RAM_R0C0_RD15), .RD14(RAM_R0C0_RD14), .RD13(RAM_R0C0_RD13), 
        .RD12(RAM_R0C0_RD12), .RD11(QX_TEMPR0_11_net), .RD10(
        QX_TEMPR0_10_net), .RD9(QX_TEMPR0_9_net), .RD8(QX_TEMPR0_8_net)
        , .RD7(QX_TEMPR0_7_net), .RD6(QX_TEMPR0_6_net), .RD5(
        QX_TEMPR0_5_net), .RD4(QX_TEMPR0_4_net), .RD3(QX_TEMPR0_3_net), 
        .RD2(QX_TEMPR0_2_net), .RD1(QX_TEMPR0_1_net), .RD0(
        QX_TEMPR0_0_net));
    OR2 ORB_GATE_10_inst (.A(ENABLE_ADDRB_10_net), .B(WEBP), .Y(
        BLKB_EN_10_net));
    AND2A AND2A_7 (.A(addr[8]), .B(addr[9]), .Y(AND2A_7_Y));
    MX2 MX2_44 (.A(MX2_16_Y), .B(MX2_86_Y), .S(BUFF_10_Y), .Y(MX2_44_Y)
        );
    MX2 MX2_56 (.A(QX_TEMPR10_1_net), .B(QX_TEMPR11_1_net), .S(
        BUFF_2_Y), .Y(MX2_56_Y));
    MX2 MX2_136 (.A(MX2_160_Y), .B(MX2_106_Y), .S(BUFF_8_Y), .Y(
        MX2_136_Y));
    NAND2 NAND2_ENABLE_ADDRB_8_inst (.A(NOR2_0_Y), .B(AND2A_5_Y), .Y(
        ENABLE_ADDRB_8_net));
    NAND2 NAND2_ENABLE_ADDRA_5_inst (.A(AND2A_2_Y), .B(AND2A_0_Y), .Y(
        ENABLE_ADDRA_5_net));
    MX2 MX2_RD_1_inst_inst_1 (.A(MX2_130_Y), .B(MX2_139_Y), .S(
        BUFF_0_Y), .Y(MX2_RD_1_inst));
    MX2 MX2_163 (.A(MX2_88_Y), .B(MX2_1_Y), .S(BUFF_8_Y), .Y(MX2_163_Y)
        );
    RAM512X18 #( .MEMORYFILE("RAM_R12C0.mem") )  RAM_R12C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_12_net), .WEN(BLKA_EN_12_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R12C0_RD17), .RD16(RAM_R12C0_RD16), .RD15(
        RAM_R12C0_RD15), .RD14(RAM_R12C0_RD14), .RD13(RAM_R12C0_RD13), 
        .RD12(RAM_R12C0_RD12), .RD11(QX_TEMPR12_11_net), .RD10(
        QX_TEMPR12_10_net), .RD9(QX_TEMPR12_9_net), .RD8(
        QX_TEMPR12_8_net), .RD7(QX_TEMPR12_7_net), .RD6(
        QX_TEMPR12_6_net), .RD5(QX_TEMPR12_5_net), .RD4(
        QX_TEMPR12_4_net), .RD3(QX_TEMPR12_3_net), .RD2(
        QX_TEMPR12_2_net), .RD1(QX_TEMPR12_1_net), .RD0(
        QX_TEMPR12_0_net));
    AND2 AND2_1 (.A(addr_0[11]), .B(addr_0[10]), .Y(AND2_1_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R4C0.mem") )  RAM_R4C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_4_net), .WEN(BLKA_EN_4_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R4C0_RD17), .RD16(RAM_R4C0_RD16), .RD15(
        RAM_R4C0_RD15), .RD14(RAM_R4C0_RD14), .RD13(RAM_R4C0_RD13), 
        .RD12(RAM_R4C0_RD12), .RD11(QX_TEMPR4_11_net), .RD10(
        QX_TEMPR4_10_net), .RD9(QX_TEMPR4_9_net), .RD8(QX_TEMPR4_8_net)
        , .RD7(QX_TEMPR4_7_net), .RD6(QX_TEMPR4_6_net), .RD5(
        QX_TEMPR4_5_net), .RD4(QX_TEMPR4_4_net), .RD3(QX_TEMPR4_3_net), 
        .RD2(QX_TEMPR4_2_net), .RD1(QX_TEMPR4_1_net), .RD0(
        QX_TEMPR4_0_net));
    AND2A AND2A_1 (.A(addr_0[10]), .B(addr_0[11]), .Y(AND2A_1_Y));
    MX2 MX2_5 (.A(MX2_164_Y), .B(MX2_79_Y), .S(BUFF_5_Y), .Y(MX2_5_Y));
    OR2 ORB_GATE_4_inst (.A(ENABLE_ADDRB_4_net), .B(WEBP), .Y(
        BLKB_EN_4_net));
    NAND2 NAND2_ENABLE_ADDRA_3_inst (.A(AND2_2_Y), .B(NOR2_1_Y), .Y(
        ENABLE_ADDRA_3_net));
    MX2 MX2_53 (.A(QX_TEMPR12_2_net), .B(QX_TEMPR13_2_net), .S(
        BUFF_13_Y), .Y(MX2_53_Y));
    MX2 MX2_25 (.A(QX_TEMPR2_5_net), .B(QX_TEMPR3_5_net), .S(BUFF_14_Y)
        , .Y(MX2_25_Y));
    MX2 MX2_161 (.A(MX2_155_Y), .B(MX2_115_Y), .S(BUFF_3_Y), .Y(
        MX2_161_Y));
    AND2A AND2A_5 (.A(addr[10]), .B(addr[11]), .Y(AND2A_5_Y));
    MX2 MX2_133 (.A(QX_TEMPR12_3_net), .B(QX_TEMPR13_3_net), .S(
        BUFF_13_Y), .Y(MX2_133_Y));
    BUFF BUFF_2 (.A(ADDRB_FF2_0_net), .Y(BUFF_2_Y));
    MX2 MX2_148 (.A(MX2_64_Y), .B(MX2_114_Y), .S(BUFF_3_Y), .Y(
        MX2_148_Y));
    NAND2 NAND2_ENABLE_ADDRA_6_inst (.A(AND2A_4_Y), .B(AND2A_0_Y), .Y(
        ENABLE_ADDRA_6_net));
    NAND2 NAND2_ENABLE_ADDRA_1_inst (.A(AND2A_2_Y), .B(NOR2_1_Y), .Y(
        ENABLE_ADDRA_1_net));
    NAND2 NAND2_ENABLE_ADDRA_15_inst (.A(AND2_2_Y), .B(AND2_1_Y), .Y(
        ENABLE_ADDRA_15_net));
    MX2 MX2_115 (.A(QX_TEMPR10_0_net), .B(QX_TEMPR11_0_net), .S(
        BUFF_11_Y), .Y(MX2_115_Y));
    MX2 MX2_61 (.A(MX2_55_Y), .B(MX2_43_Y), .S(BUFF_16_Y), .Y(MX2_61_Y)
        );
    MX2 MX2_147 (.A(MX2_0_Y), .B(MX2_159_Y), .S(BUFF_8_Y), .Y(
        MX2_147_Y));
    MX2 MX2_82 (.A(QX_TEMPR14_0_net), .B(QX_TEMPR15_0_net), .S(
        BUFF_11_Y), .Y(MX2_82_Y));
    MX2 MX2_131 (.A(QX_TEMPR4_7_net), .B(QX_TEMPR5_7_net), .S(BUFF_4_Y)
        , .Y(MX2_131_Y));
    NAND2 NAND2_ENABLE_ADDRA_4_inst (.A(NOR2_2_Y), .B(AND2A_0_Y), .Y(
        ENABLE_ADDRA_4_net));
    NOR2 NOR2_3 (.A(addr[11]), .B(addr[10]), .Y(NOR2_3_Y));
    OR2 ORA_GATE_4_inst (.A(ENABLE_ADDRA_4_net), .B(WEAP), .Y(
        BLKA_EN_4_net));
    MX2 MX2_57 (.A(QX_TEMPR6_11_net), .B(QX_TEMPR7_11_net), .S(
        BUFF_7_Y), .Y(MX2_57_Y));
    MX2 MX2_71 (.A(QX_TEMPR10_8_net), .B(QX_TEMPR11_8_net), .S(
        BUFF_1_Y), .Y(MX2_71_Y));
    INV WEBUBBLEB (.A(top_code_0_n_rd_en), .Y(WEBP));
    MX2 MX2_20 (.A(QX_TEMPR0_4_net), .B(QX_TEMPR1_4_net), .S(BUFF_13_Y)
        , .Y(MX2_20_Y));
    MX2 MX2_19 (.A(QX_TEMPR4_3_net), .B(QX_TEMPR5_3_net), .S(BUFF_13_Y)
        , .Y(MX2_19_Y));
    OR2 ORA_GATE_13_inst (.A(ENABLE_ADDRA_13_net), .B(WEAP), .Y(
        BLKA_EN_13_net));
    NAND2 NAND2_ENABLE_ADDRA_13_inst (.A(AND2A_2_Y), .B(AND2_1_Y), .Y(
        ENABLE_ADDRA_13_net));
    OR2 ORB_GATE_5_inst (.A(ENABLE_ADDRB_5_net), .B(WEBP), .Y(
        BLKB_EN_5_net));
    MX2 MX2_88 (.A(QX_TEMPR8_6_net), .B(QX_TEMPR9_6_net), .S(BUFF_12_Y)
        , .Y(MX2_88_Y));
    MX2 MX2_31 (.A(QX_TEMPR14_1_net), .B(QX_TEMPR15_1_net), .S(
        BUFF_2_Y), .Y(MX2_31_Y));
    OR2 ORB_GATE_2_inst (.A(ENABLE_ADDRB_2_net), .B(WEBP), .Y(
        BLKB_EN_2_net));
    MX2 MX2_155 (.A(QX_TEMPR8_0_net), .B(QX_TEMPR9_0_net), .S(
        BUFF_11_Y), .Y(MX2_155_Y));
    MX2 MX2_14 (.A(MX2_110_Y), .B(MX2_25_Y), .S(BUFF_8_Y), .Y(MX2_14_Y)
        );
    MX2 MX2_65 (.A(MX2_90_Y), .B(MX2_38_Y), .S(BUFF_18_Y), .Y(MX2_65_Y)
        );
    NAND2 NAND2_ENABLE_ADDRB_10_inst (.A(AND2A_7_Y), .B(AND2A_5_Y), .Y(
        ENABLE_ADDRB_10_net));
    GND GND_i (.Y(GND));
    MX2 MX2_91 (.A(MX2_156_Y), .B(MX2_54_Y), .S(BUFF_18_Y), .Y(
        MX2_91_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R9C0.mem") )  RAM_R9C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_9_net), .WEN(BLKA_EN_9_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R9C0_RD17), .RD16(RAM_R9C0_RD16), .RD15(
        RAM_R9C0_RD15), .RD14(RAM_R9C0_RD14), .RD13(RAM_R9C0_RD13), 
        .RD12(RAM_R9C0_RD12), .RD11(QX_TEMPR9_11_net), .RD10(
        QX_TEMPR9_10_net), .RD9(QX_TEMPR9_9_net), .RD8(QX_TEMPR9_8_net)
        , .RD7(QX_TEMPR9_7_net), .RD6(QX_TEMPR9_6_net), .RD5(
        QX_TEMPR9_5_net), .RD4(QX_TEMPR9_4_net), .RD3(QX_TEMPR9_3_net), 
        .RD2(QX_TEMPR9_2_net), .RD1(QX_TEMPR9_1_net), .RD0(
        QX_TEMPR9_0_net));
    MX2 MX2_75 (.A(QX_TEMPR0_3_net), .B(QX_TEMPR1_3_net), .S(BUFF_13_Y)
        , .Y(MX2_75_Y));
    MX2 MX2_86 (.A(MX2_23_Y), .B(MX2_126_Y), .S(BUFF_5_Y), .Y(MX2_86_Y)
        );
    BUFF BUFF_14 (.A(ADDRB_FF2_0_net), .Y(BUFF_14_Y));
    OR2 ORB_GATE_9_inst (.A(ENABLE_ADDRB_9_net), .B(WEBP), .Y(
        BLKB_EN_9_net));
    VCC VCC_i_0 (.Y(VCC_0));
    MX2 MX2_142 (.A(MX2_49_Y), .B(MX2_10_Y), .S(BUFF_3_Y), .Y(
        MX2_142_Y));
    OR2 ORA_GATE_5_inst (.A(ENABLE_ADDRA_5_net), .B(WEAP), .Y(
        BLKA_EN_5_net));
    NOR2 NOR2_0 (.A(addr[9]), .B(addr[8]), .Y(NOR2_0_Y));
    OR2 ORB_GATE_1_inst (.A(ENABLE_ADDRB_1_net), .B(WEBP), .Y(
        BLKB_EN_1_net));
    OR2 ORB_GATE_12_inst (.A(ENABLE_ADDRB_12_net), .B(WEBP), .Y(
        BLKB_EN_12_net));
    MX2 MX2_35 (.A(MX2_26_Y), .B(MX2_109_Y), .S(BUFF_15_Y), .Y(
        MX2_35_Y));
    OR2 ORA_GATE_2_inst (.A(ENABLE_ADDRA_2_net), .B(WEAP), .Y(
        BLKA_EN_2_net));
    MX2 MX2_8 (.A(QX_TEMPR14_2_net), .B(QX_TEMPR15_2_net), .S(
        BUFF_13_Y), .Y(MX2_8_Y));
    MX2 MX2_105 (.A(MX2_123_Y), .B(MX2_74_Y), .S(BUFF_5_Y), .Y(
        MX2_105_Y));
    MX2 MX2_60 (.A(QX_TEMPR10_7_net), .B(QX_TEMPR11_7_net), .S(
        BUFF_4_Y), .Y(MX2_60_Y));
    MX2 MX2_83 (.A(QX_TEMPR12_7_net), .B(QX_TEMPR13_7_net), .S(
        BUFF_4_Y), .Y(MX2_83_Y));
    MX2 MX2_RD_0_inst_inst_1 (.A(MX2_165_Y), .B(MX2_34_Y), .S(BUFF_0_Y)
        , .Y(MX2_RD_0_inst));
    MX2 MX2_RD_4_inst_inst_1 (.A(MX2_89_Y), .B(MX2_87_Y), .S(BUFF_0_Y), 
        .Y(MX2_RD_4_inst));
    MX2 MX2_114 (.A(QX_TEMPR2_0_net), .B(QX_TEMPR3_0_net), .S(
        BUFF_11_Y), .Y(MX2_114_Y));
    MX2 MX2_RD_8_inst_inst_1 (.A(MX2_30_Y), .B(MX2_152_Y), .S(BUFF_9_Y)
        , .Y(MX2_RD_8_inst));
    MX2 MX2_110 (.A(QX_TEMPR0_5_net), .B(QX_TEMPR1_5_net), .S(
        BUFF_14_Y), .Y(MX2_110_Y));
    MX2 MX2_95 (.A(QX_TEMPR2_7_net), .B(QX_TEMPR3_7_net), .S(BUFF_4_Y), 
        .Y(MX2_95_Y));
    MX2 MX2_119 (.A(QX_TEMPR4_11_net), .B(QX_TEMPR5_11_net), .S(
        BUFF_7_Y), .Y(MX2_119_Y));
    AND2 AND2_3 (.A(addr[11]), .B(addr[10]), .Y(AND2_3_Y));
    MX2 MX2_70 (.A(QX_TEMPR6_9_net), .B(QX_TEMPR7_9_net), .S(BUFF_1_Y), 
        .Y(MX2_70_Y));
    OR2 ORA_GATE_9_inst (.A(ENABLE_ADDRA_9_net), .B(WEAP), .Y(
        BLKA_EN_9_net));
    NAND2 NAND2_ENABLE_ADDRA_12_inst (.A(NOR2_2_Y), .B(AND2_1_Y), .Y(
        ENABLE_ADDRA_12_net));
    NAND2 NAND2_ENABLE_ADDRA_14_inst (.A(AND2A_4_Y), .B(AND2_1_Y), .Y(
        ENABLE_ADDRA_14_net));
    MX2 MX2_146 (.A(QX_TEMPR4_0_net), .B(QX_TEMPR5_0_net), .S(
        BUFF_11_Y), .Y(MX2_146_Y));
    MX2 MX2_59 (.A(QX_TEMPR0_8_net), .B(QX_TEMPR1_8_net), .S(BUFF_4_Y), 
        .Y(MX2_59_Y));
    OR2 ORA_GATE_1_inst (.A(ENABLE_ADDRA_1_net), .B(WEAP), .Y(
        BLKA_EN_1_net));
    BUFF BUFF_5 (.A(ADDRB_FF2_1_net), .Y(BUFF_5_Y));
    MX2 MX2_30 (.A(MX2_103_Y), .B(MX2_91_Y), .S(BUFF_10_Y), .Y(
        MX2_30_Y));
    MX2 MX2_22 (.A(QX_TEMPR8_9_net), .B(QX_TEMPR9_9_net), .S(BUFF_6_Y), 
        .Y(MX2_22_Y));
    OR2 ORB_GATE_6_inst (.A(ENABLE_ADDRB_6_net), .B(WEBP), .Y(
        BLKB_EN_6_net));
    MX2 MX2_87 (.A(MX2_124_Y), .B(MX2_2_Y), .S(BUFF_17_Y), .Y(MX2_87_Y)
        );
    VCC VCC_i (.Y(VCC));
    MX2 MX2_154 (.A(MX2_158_Y), .B(MX2_9_Y), .S(BUFF_10_Y), .Y(
        MX2_154_Y));
    NOR2 NOR2_1 (.A(addr_0[11]), .B(addr_0[10]), .Y(NOR2_1_Y));
    MX2 MX2_90 (.A(QX_TEMPR12_8_net), .B(QX_TEMPR13_8_net), .S(
        BUFF_1_Y), .Y(MX2_90_Y));
    MX2 MX2_54 (.A(QX_TEMPR6_8_net), .B(QX_TEMPR7_8_net), .S(BUFF_1_Y), 
        .Y(MX2_54_Y));
    MX2 MX2_150 (.A(QX_TEMPR0_7_net), .B(QX_TEMPR1_7_net), .S(BUFF_4_Y)
        , .Y(MX2_150_Y));
    MX2 MX2_159 (.A(QX_TEMPR6_5_net), .B(QX_TEMPR7_5_net), .S(
        BUFF_14_Y), .Y(MX2_159_Y));
    NAND2 NAND2_ENABLE_ADDRA_7_inst (.A(AND2_2_Y), .B(AND2A_0_Y), .Y(
        ENABLE_ADDRA_7_net));
    MX2 MX2_0 (.A(QX_TEMPR4_5_net), .B(QX_TEMPR5_5_net), .S(BUFF_14_Y), 
        .Y(MX2_0_Y));
    MX2 MX2_143 (.A(MX2_76_Y), .B(MX2_51_Y), .S(BUFF_17_Y), .Y(
        MX2_143_Y));
    DFN1 BFF1_1_inst (.D(addr[9]), .CLK(n_rdclk), .Q(ADDRB_FF2_1_net));
    NAND2 NAND2_ENABLE_ADDRB_7_inst (.A(AND2_0_Y), .B(AND2A_3_Y), .Y(
        ENABLE_ADDRB_7_net));
    MX2 MX2_41 (.A(QX_TEMPR10_11_net), .B(QX_TEMPR11_11_net), .S(
        BUFF_7_Y), .Y(MX2_41_Y));
    MX2 MX2_28 (.A(MX2_18_Y), .B(MX2_96_Y), .S(BUFF_5_Y), .Y(MX2_28_Y));
    OR2 ORA_GATE_6_inst (.A(ENABLE_ADDRA_6_net), .B(WEAP), .Y(
        BLKA_EN_6_net));
    MX2 MX2_141 (.A(QX_TEMPR6_2_net), .B(QX_TEMPR7_2_net), .S(BUFF_2_Y)
        , .Y(MX2_141_Y));
    NAND2 NAND2_ENABLE_ADDRB_4_inst (.A(NOR2_0_Y), .B(AND2A_3_Y), .Y(
        ENABLE_ADDRB_4_net));
    MX2 MX2_104 (.A(QX_TEMPR2_9_net), .B(QX_TEMPR3_9_net), .S(BUFF_1_Y)
        , .Y(MX2_104_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R2C0.mem") )  RAM_R2C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_2_net), .WEN(BLKA_EN_2_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R2C0_RD17), .RD16(RAM_R2C0_RD16), .RD15(
        RAM_R2C0_RD15), .RD14(RAM_R2C0_RD14), .RD13(RAM_R2C0_RD13), 
        .RD12(RAM_R2C0_RD12), .RD11(QX_TEMPR2_11_net), .RD10(
        QX_TEMPR2_10_net), .RD9(QX_TEMPR2_9_net), .RD8(QX_TEMPR2_8_net)
        , .RD7(QX_TEMPR2_7_net), .RD6(QX_TEMPR2_6_net), .RD5(
        QX_TEMPR2_5_net), .RD4(QX_TEMPR2_4_net), .RD3(QX_TEMPR2_3_net), 
        .RD2(QX_TEMPR2_2_net), .RD1(QX_TEMPR2_1_net), .RD0(
        QX_TEMPR2_0_net));
    MX2 MX2_100 (.A(QX_TEMPR6_0_net), .B(QX_TEMPR7_0_net), .S(
        BUFF_11_Y), .Y(MX2_100_Y));
    MX2 MX2_26 (.A(MX2_62_Y), .B(MX2_117_Y), .S(BUFF_16_Y), .Y(
        MX2_26_Y));
    MX2 MX2_109 (.A(MX2_133_Y), .B(MX2_85_Y), .S(BUFF_16_Y), .Y(
        MX2_109_Y));
    AND2A AND2A_2 (.A(addr_0[9]), .B(addr_0[8]), .Y(AND2A_2_Y));
    MX2 MX2_125 (.A(QX_TEMPR4_4_net), .B(QX_TEMPR5_4_net), .S(
        BUFF_14_Y), .Y(MX2_125_Y));
    MX2 MX2_62 (.A(QX_TEMPR8_3_net), .B(QX_TEMPR9_3_net), .S(BUFF_13_Y)
        , .Y(MX2_62_Y));
    MX2 MX2_45 (.A(QX_TEMPR8_1_net), .B(QX_TEMPR9_1_net), .S(BUFF_2_Y), 
        .Y(MX2_45_Y));
    MX2 MX2_118 (.A(MX2_61_Y), .B(MX2_39_Y), .S(BUFF_15_Y), .Y(
        MX2_118_Y));
    MX2 MX2_2 (.A(MX2_29_Y), .B(MX2_134_Y), .S(BUFF_16_Y), .Y(MX2_2_Y));
    MX2 MX2_72 (.A(QX_TEMPR6_7_net), .B(QX_TEMPR7_7_net), .S(BUFF_4_Y), 
        .Y(MX2_72_Y));
    NAND2 NAND2_ENABLE_ADDRB_15_inst (.A(AND2_0_Y), .B(AND2_3_Y), .Y(
        ENABLE_ADDRB_15_net));
    MX2 MX2_RD_10_inst_inst_1 (.A(MX2_44_Y), .B(MX2_81_Y), .S(BUFF_9_Y)
        , .Y(MX2_RD_10_inst));
    MX2 MX2_23 (.A(QX_TEMPR4_10_net), .B(QX_TEMPR5_10_net), .S(
        BUFF_6_Y), .Y(MX2_23_Y));
    NAND2 NAND2_ENABLE_ADDRB_6_inst (.A(AND2A_7_Y), .B(AND2A_3_Y), .Y(
        ENABLE_ADDRB_6_net));
    MX2 MX2_117 (.A(QX_TEMPR10_3_net), .B(QX_TEMPR11_3_net), .S(
        BUFF_13_Y), .Y(MX2_117_Y));
    OR2 ORB_GATE_7_inst (.A(ENABLE_ADDRB_7_net), .B(WEBP), .Y(
        BLKB_EN_7_net));
    BUFF BUFF_12 (.A(ADDRB_FF2_0_net), .Y(BUFF_12_Y));
    AND2A AND2A_4 (.A(addr_0[8]), .B(addr_0[9]), .Y(AND2A_4_Y));
    MX2 MX2_68 (.A(MX2_149_Y), .B(MX2_138_Y), .S(BUFF_15_Y), .Y(
        MX2_68_Y));
    MX2 MX2_RD_3_inst_inst_1 (.A(MX2_68_Y), .B(MX2_35_Y), .S(BUFF_0_Y), 
        .Y(MX2_RD_3_inst));
    MX2 MX2_32 (.A(MX2_162_Y), .B(MX2_105_Y), .S(BUFF_10_Y), .Y(
        MX2_32_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R14C0.mem") )  RAM_R14C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_14_net), .WEN(BLKA_EN_14_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R14C0_RD17), .RD16(RAM_R14C0_RD16), .RD15(
        RAM_R14C0_RD15), .RD14(RAM_R14C0_RD14), .RD13(RAM_R14C0_RD13), 
        .RD12(RAM_R14C0_RD12), .RD11(QX_TEMPR14_11_net), .RD10(
        QX_TEMPR14_10_net), .RD9(QX_TEMPR14_9_net), .RD8(
        QX_TEMPR14_8_net), .RD7(QX_TEMPR14_7_net), .RD6(
        QX_TEMPR14_6_net), .RD5(QX_TEMPR14_5_net), .RD4(
        QX_TEMPR14_4_net), .RD3(QX_TEMPR14_3_net), .RD2(
        QX_TEMPR14_2_net), .RD1(QX_TEMPR14_1_net), .RD0(
        QX_TEMPR14_0_net));
    MX2 MX2_89 (.A(MX2_40_Y), .B(MX2_92_Y), .S(BUFF_17_Y), .Y(MX2_89_Y)
        );
    OR2 ORB_GATE_15_inst (.A(ENABLE_ADDRB_15_net), .B(WEBP), .Y(
        BLKB_EN_15_net));
    NAND2 NAND2_ENABLE_ADDRB_13_inst (.A(AND2A_6_Y), .B(AND2_3_Y), .Y(
        ENABLE_ADDRB_13_net));
    MX2 MX2_RD_2_inst_inst_1 (.A(MX2_122_Y), .B(MX2_118_Y), .S(
        BUFF_0_Y), .Y(MX2_RD_2_inst));
    OR2 ORB_GATE_8_inst (.A(ENABLE_ADDRB_8_net), .B(WEBP), .Y(
        BLKB_EN_8_net));
    MX2 MX2_78 (.A(QX_TEMPR12_1_net), .B(QX_TEMPR13_1_net), .S(
        BUFF_2_Y), .Y(MX2_78_Y));
    BUFF BUFF_0 (.A(ADDRB_FF2_3_net), .Y(BUFF_0_Y));
    MX2 MX2_40 (.A(MX2_20_Y), .B(MX2_52_Y), .S(BUFF_16_Y), .Y(MX2_40_Y)
        );
    RAM512X18 #( .MEMORYFILE("RAM_R8C0.mem") )  RAM_R8C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_8_net), .WEN(BLKA_EN_8_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R8C0_RD17), .RD16(RAM_R8C0_RD16), .RD15(
        RAM_R8C0_RD15), .RD14(RAM_R8C0_RD14), .RD13(RAM_R8C0_RD13), 
        .RD12(RAM_R8C0_RD12), .RD11(QX_TEMPR8_11_net), .RD10(
        QX_TEMPR8_10_net), .RD9(QX_TEMPR8_9_net), .RD8(QX_TEMPR8_8_net)
        , .RD7(QX_TEMPR8_7_net), .RD6(QX_TEMPR8_6_net), .RD5(
        QX_TEMPR8_5_net), .RD4(QX_TEMPR8_4_net), .RD3(QX_TEMPR8_3_net), 
        .RD2(QX_TEMPR8_2_net), .RD1(QX_TEMPR8_1_net), .RD0(
        QX_TEMPR8_0_net));
    MX2 MX2_92 (.A(MX2_125_Y), .B(MX2_63_Y), .S(BUFF_16_Y), .Y(
        MX2_92_Y));
    MX2 MX2_158 (.A(MX2_80_Y), .B(MX2_166_Y), .S(BUFF_5_Y), .Y(
        MX2_158_Y));
    INV WEBUBBLEA (.A(n_acq_change_0_n_acq_start), .Y(WEAP));
    MX2 MX2_27 (.A(MX2_131_Y), .B(MX2_72_Y), .S(BUFF_8_Y), .Y(MX2_27_Y)
        );
    MX2 MX2_165 (.A(MX2_148_Y), .B(MX2_6_Y), .S(BUFF_15_Y), .Y(
        MX2_165_Y));
    MX2 MX2_66 (.A(MX2_36_Y), .B(MX2_107_Y), .S(BUFF_17_Y), .Y(
        MX2_66_Y));
    MX2 MX2_84 (.A(MX2_45_Y), .B(MX2_56_Y), .S(BUFF_3_Y), .Y(MX2_84_Y));
    MX2 MX2_11 (.A(MX2_93_Y), .B(MX2_41_Y), .S(BUFF_5_Y), .Y(MX2_11_Y));
    OR2 ORA_GATE_15_inst (.A(ENABLE_ADDRA_15_net), .B(WEAP), .Y(
        BLKA_EN_15_net));
    MX2 MX2_157 (.A(MX2_24_Y), .B(MX2_121_Y), .S(BUFF_8_Y), .Y(
        MX2_157_Y));
    OR2 ORA_GATE_7_inst (.A(ENABLE_ADDRA_7_net), .B(WEAP), .Y(
        BLKA_EN_7_net));
    MX2 MX2_38 (.A(QX_TEMPR14_8_net), .B(QX_TEMPR15_8_net), .S(
        BUFF_1_Y), .Y(MX2_38_Y));
    MX2 MX2_76 (.A(MX2_101_Y), .B(MX2_60_Y), .S(BUFF_18_Y), .Y(
        MX2_76_Y));
    MX2 MX2_6 (.A(MX2_146_Y), .B(MX2_100_Y), .S(BUFF_3_Y), .Y(MX2_6_Y));
    MX2 MX2_135 (.A(MX2_128_Y), .B(MX2_47_Y), .S(BUFF_5_Y), .Y(
        MX2_135_Y));
    MX2 MX2_112 (.A(QX_TEMPR6_6_net), .B(QX_TEMPR7_6_net), .S(
        BUFF_12_Y), .Y(MX2_112_Y));
    MX2 MX2_98 (.A(MX2_150_Y), .B(MX2_95_Y), .S(BUFF_8_Y), .Y(MX2_98_Y)
        );
    MX2 MX2_63 (.A(QX_TEMPR6_4_net), .B(QX_TEMPR7_4_net), .S(BUFF_14_Y)
        , .Y(MX2_63_Y));
    OR2 ORA_GATE_8_inst (.A(ENABLE_ADDRA_8_net), .B(WEAP), .Y(
        BLKA_EN_8_net));
    NAND2 NAND2_ENABLE_ADDRB_3_inst (.A(AND2_0_Y), .B(NOR2_3_Y), .Y(
        ENABLE_ADDRB_3_net));
    MX2 MX2_124 (.A(MX2_137_Y), .B(MX2_7_Y), .S(BUFF_16_Y), .Y(
        MX2_124_Y));
    OR2 ORA_GATE_11_inst (.A(ENABLE_ADDRA_11_net), .B(WEAP), .Y(
        BLKA_EN_11_net));
    MX2 MX2_36 (.A(MX2_42_Y), .B(MX2_37_Y), .S(BUFF_8_Y), .Y(MX2_36_Y));
    MX2 MX2_120 (.A(QX_TEMPR2_8_net), .B(QX_TEMPR3_8_net), .S(BUFF_4_Y)
        , .Y(MX2_120_Y));
    MX2 MX2_129 (.A(QX_TEMPR0_1_net), .B(QX_TEMPR1_1_net), .S(
        BUFF_11_Y), .Y(MX2_129_Y));
    MX2 MX2_108 (.A(MX2_132_Y), .B(MX2_82_Y), .S(BUFF_3_Y), .Y(
        MX2_108_Y));
    MX2 MX2_RD_7_inst_inst_1 (.A(MX2_116_Y), .B(MX2_143_Y), .S(
        BUFF_9_Y), .Y(MX2_RD_7_inst));
    MX2 MX2_7 (.A(QX_TEMPR10_4_net), .B(QX_TEMPR11_4_net), .S(
        BUFF_14_Y), .Y(MX2_7_Y));
    AND2A AND2A_3 (.A(addr[11]), .B(addr[10]), .Y(AND2A_3_Y));
    NAND2 NAND2_ENABLE_ADDRA_0_inst (.A(NOR2_2_Y), .B(NOR2_1_Y), .Y(
        ENABLE_ADDRA_0_net));
    MX2 MX2_73 (.A(MX2_67_Y), .B(MX2_151_Y), .S(BUFF_3_Y), .Y(MX2_73_Y)
        );
    BUFF BUFF_9 (.A(ADDRB_FF2_3_net), .Y(BUFF_9_Y));
    MX2 MX2_15 (.A(QX_TEMPR4_6_net), .B(QX_TEMPR5_6_net), .S(BUFF_12_Y)
        , .Y(MX2_15_Y));
    MX2 MX2_107 (.A(MX2_15_Y), .B(MX2_112_Y), .S(BUFF_8_Y), .Y(
        MX2_107_Y));
    AND2A AND2A_6 (.A(addr[9]), .B(addr[8]), .Y(AND2A_6_Y));
    MX2 MX2_96 (.A(QX_TEMPR14_10_net), .B(QX_TEMPR15_10_net), .S(
        BUFF_7_Y), .Y(MX2_96_Y));
    MX2 MX2_3 (.A(QX_TEMPR0_10_net), .B(QX_TEMPR1_10_net), .S(BUFF_6_Y)
        , .Y(MX2_3_Y));
    MX2 MX2_33 (.A(QX_TEMPR14_7_net), .B(QX_TEMPR15_7_net), .S(
        BUFF_4_Y), .Y(MX2_33_Y));
    OR2 ORA_GATE_14_inst (.A(ENABLE_ADDRA_14_net), .B(WEAP), .Y(
        BLKA_EN_14_net));
    MX2 MX2_67 (.A(QX_TEMPR0_2_net), .B(QX_TEMPR1_2_net), .S(BUFF_2_Y), 
        .Y(MX2_67_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R13C0.mem") )  RAM_R13C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_13_net), .WEN(BLKA_EN_13_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R13C0_RD17), .RD16(RAM_R13C0_RD16), .RD15(
        RAM_R13C0_RD15), .RD14(RAM_R13C0_RD14), .RD13(RAM_R13C0_RD13), 
        .RD12(RAM_R13C0_RD12), .RD11(QX_TEMPR13_11_net), .RD10(
        QX_TEMPR13_10_net), .RD9(QX_TEMPR13_9_net), .RD8(
        QX_TEMPR13_8_net), .RD7(QX_TEMPR13_7_net), .RD6(
        QX_TEMPR13_6_net), .RD5(QX_TEMPR13_5_net), .RD4(
        QX_TEMPR13_4_net), .RD3(QX_TEMPR13_3_net), .RD2(
        QX_TEMPR13_2_net), .RD1(QX_TEMPR13_1_net), .RD0(
        QX_TEMPR13_0_net));
    MX2 MX2_152 (.A(MX2_102_Y), .B(MX2_65_Y), .S(BUFF_10_Y), .Y(
        MX2_152_Y));
    GND GND_i_0 (.Y(GND_0));
    OR2 ORB_GATE_14_inst (.A(ENABLE_ADDRB_14_net), .B(WEBP), .Y(
        BLKB_EN_14_net));
    NAND2 NAND2_ENABLE_ADDRB_12_inst (.A(NOR2_0_Y), .B(AND2_3_Y), .Y(
        ENABLE_ADDRB_12_net));
    NAND2 NAND2_ENABLE_ADDRB_14_inst (.A(AND2A_7_Y), .B(AND2_3_Y), .Y(
        ENABLE_ADDRB_14_net));
    MX2 MX2_116 (.A(MX2_98_Y), .B(MX2_27_Y), .S(BUFF_17_Y), .Y(
        MX2_116_Y));
    BUFF BUFF_6 (.A(ADDRB_FF2_0_net), .Y(BUFF_6_Y));
    MX2 MX2_9 (.A(MX2_119_Y), .B(MX2_57_Y), .S(BUFF_5_Y), .Y(MX2_9_Y));
    BUFF BUFF_7 (.A(ADDRB_FF2_0_net), .Y(BUFF_7_Y));
    NAND2 NAND2_ENABLE_ADDRA_11_inst (.A(AND2_2_Y), .B(AND2A_1_Y), .Y(
        ENABLE_ADDRA_11_net));
    MX2 MX2_93 (.A(QX_TEMPR8_11_net), .B(QX_TEMPR9_11_net), .S(
        BUFF_7_Y), .Y(MX2_93_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R11C0.mem") )  RAM_R11C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_11_net), .WEN(BLKA_EN_11_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R11C0_RD17), .RD16(RAM_R11C0_RD16), .RD15(
        RAM_R11C0_RD15), .RD14(RAM_R11C0_RD14), .RD13(RAM_R11C0_RD13), 
        .RD12(RAM_R11C0_RD12), .RD11(QX_TEMPR11_11_net), .RD10(
        QX_TEMPR11_10_net), .RD9(QX_TEMPR11_9_net), .RD8(
        QX_TEMPR11_8_net), .RD7(QX_TEMPR11_7_net), .RD6(
        QX_TEMPR11_6_net), .RD5(QX_TEMPR11_5_net), .RD4(
        QX_TEMPR11_4_net), .RD3(QX_TEMPR11_3_net), .RD2(
        QX_TEMPR11_2_net), .RD1(QX_TEMPR11_1_net), .RD0(
        QX_TEMPR11_0_net));
    MX2 MX2_77 (.A(MX2_163_Y), .B(MX2_157_Y), .S(BUFF_17_Y), .Y(
        MX2_77_Y));
    AND2A AND2A_0 (.A(addr_0[11]), .B(addr_0[10]), .Y(AND2A_0_Y));
    BUFF BUFF_16 (.A(ADDRB_FF2_1_net), .Y(BUFF_16_Y));
    MX2 MX2_10 (.A(QX_TEMPR6_1_net), .B(QX_TEMPR7_1_net), .S(BUFF_2_Y), 
        .Y(MX2_10_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R15C0.mem") )  RAM_R15C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_15_net), .WEN(BLKA_EN_15_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R15C0_RD17), .RD16(RAM_R15C0_RD16), .RD15(
        RAM_R15C0_RD15), .RD14(RAM_R15C0_RD14), .RD13(RAM_R15C0_RD13), 
        .RD12(RAM_R15C0_RD12), .RD11(QX_TEMPR15_11_net), .RD10(
        QX_TEMPR15_10_net), .RD9(QX_TEMPR15_9_net), .RD8(
        QX_TEMPR15_8_net), .RD7(QX_TEMPR15_7_net), .RD6(
        QX_TEMPR15_6_net), .RD5(QX_TEMPR15_5_net), .RD4(
        QX_TEMPR15_4_net), .RD3(QX_TEMPR15_3_net), .RD2(
        QX_TEMPR15_2_net), .RD1(QX_TEMPR15_1_net), .RD0(
        QX_TEMPR15_0_net));
    MX2 MX2_164 (.A(QX_TEMPR12_11_net), .B(QX_TEMPR13_11_net), .S(
        BUFF_7_Y), .Y(MX2_164_Y));
    MX2 MX2_160 (.A(QX_TEMPR12_5_net), .B(QX_TEMPR13_5_net), .S(
        BUFF_12_Y), .Y(MX2_160_Y));
    BUFF BUFF_17 (.A(ADDRB_FF2_2_net), .Y(BUFF_17_Y));
    NAND2 NAND2_ENABLE_ADDRA_2_inst (.A(AND2A_4_Y), .B(NOR2_1_Y), .Y(
        ENABLE_ADDRA_2_net));
    MX2 MX2_42 (.A(QX_TEMPR0_6_net), .B(QX_TEMPR1_6_net), .S(BUFF_12_Y)
        , .Y(MX2_42_Y));
    MX2 MX2_51 (.A(MX2_83_Y), .B(MX2_33_Y), .S(BUFF_18_Y), .Y(MX2_51_Y)
        );
    MX2 MX2_29 (.A(QX_TEMPR12_4_net), .B(QX_TEMPR13_4_net), .S(
        BUFF_14_Y), .Y(MX2_29_Y));
    MX2 MX2_RD_6_inst_inst_1 (.A(MX2_66_Y), .B(MX2_77_Y), .S(BUFF_9_Y), 
        .Y(MX2_RD_6_inst));
    MX2 MX2_37 (.A(QX_TEMPR2_6_net), .B(QX_TEMPR3_6_net), .S(BUFF_12_Y)
        , .Y(MX2_37_Y));
    MX2 MX2_113 (.A(MX2_12_Y), .B(MX2_144_Y), .S(BUFF_8_Y), .Y(
        MX2_113_Y));
    MX2 MX2_102 (.A(MX2_13_Y), .B(MX2_71_Y), .S(BUFF_18_Y), .Y(
        MX2_102_Y));
    AND2 AND2_0 (.A(addr[9]), .B(addr[8]), .Y(AND2_0_Y));
    MX2 MX2_156 (.A(QX_TEMPR4_8_net), .B(QX_TEMPR5_8_net), .S(BUFF_1_Y)
        , .Y(MX2_156_Y));
    MX2 MX2_134 (.A(QX_TEMPR14_4_net), .B(QX_TEMPR15_4_net), .S(
        BUFF_14_Y), .Y(MX2_134_Y));
    BUFF BUFF_3 (.A(ADDRB_FF2_1_net), .Y(BUFF_3_Y));
    MX2 MX2_97 (.A(MX2_153_Y), .B(MX2_70_Y), .S(BUFF_18_Y), .Y(
        MX2_97_Y));
    MX2 MX2_130 (.A(MX2_94_Y), .B(MX2_142_Y), .S(BUFF_15_Y), .Y(
        MX2_130_Y));
    MX2 MX2_24 (.A(QX_TEMPR12_6_net), .B(QX_TEMPR13_6_net), .S(
        BUFF_12_Y), .Y(MX2_24_Y));
    MX2 MX2_139 (.A(MX2_84_Y), .B(MX2_46_Y), .S(BUFF_15_Y), .Y(
        MX2_139_Y));
    MX2 MX2_111 (.A(QX_TEMPR10_9_net), .B(QX_TEMPR11_9_net), .S(
        BUFF_6_Y), .Y(MX2_111_Y));
    OR2 ORA_GATE_12_inst (.A(ENABLE_ADDRA_12_net), .B(WEAP), .Y(
        BLKA_EN_12_net));
    MX2 MX2_48 (.A(MX2_113_Y), .B(MX2_136_Y), .S(BUFF_17_Y), .Y(
        MX2_48_Y));
    DFN1 BFF1_0_inst (.D(addr[8]), .CLK(n_rdclk), .Q(ADDRB_FF2_0_net));
    RAM512X18 #( .MEMORYFILE("RAM_R1C0.mem") )  RAM_R1C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_1_net), .WEN(BLKA_EN_1_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R1C0_RD17), .RD16(RAM_R1C0_RD16), .RD15(
        RAM_R1C0_RD15), .RD14(RAM_R1C0_RD14), .RD13(RAM_R1C0_RD13), 
        .RD12(RAM_R1C0_RD12), .RD11(QX_TEMPR1_11_net), .RD10(
        QX_TEMPR1_10_net), .RD9(QX_TEMPR1_9_net), .RD8(QX_TEMPR1_8_net)
        , .RD7(QX_TEMPR1_7_net), .RD6(QX_TEMPR1_6_net), .RD5(
        QX_TEMPR1_5_net), .RD4(QX_TEMPR1_4_net), .RD3(QX_TEMPR1_3_net), 
        .RD2(QX_TEMPR1_2_net), .RD1(QX_TEMPR1_1_net), .RD0(
        QX_TEMPR1_0_net));
    MX2 MX2_55 (.A(QX_TEMPR8_2_net), .B(QX_TEMPR9_2_net), .S(BUFF_2_Y), 
        .Y(MX2_55_Y));
    MX2 MX2_128 (.A(QX_TEMPR8_10_net), .B(QX_TEMPR9_10_net), .S(
        BUFF_6_Y), .Y(MX2_128_Y));
    MX2 MX2_153 (.A(QX_TEMPR4_9_net), .B(QX_TEMPR5_9_net), .S(BUFF_1_Y)
        , .Y(MX2_153_Y));
    MX2 MX2_127 (.A(QX_TEMPR2_3_net), .B(QX_TEMPR3_3_net), .S(
        BUFF_13_Y), .Y(MX2_127_Y));
    MX2 MX2_46 (.A(MX2_78_Y), .B(MX2_31_Y), .S(BUFF_3_Y), .Y(MX2_46_Y));
    MX2 MX2_106 (.A(QX_TEMPR14_5_net), .B(QX_TEMPR15_5_net), .S(
        BUFF_12_Y), .Y(MX2_106_Y));
    MX2 MX2_RD_5_inst_inst_1 (.A(MX2_140_Y), .B(MX2_48_Y), .S(BUFF_0_Y)
        , .Y(MX2_RD_5_inst));
    MX2 MX2_RD_9_inst_inst_1 (.A(MX2_50_Y), .B(MX2_32_Y), .S(BUFF_9_Y), 
        .Y(MX2_RD_9_inst));
    BUFF BUFF_15 (.A(ADDRB_FF2_2_net), .Y(BUFF_15_Y));
    MX2 MX2_69 (.A(QX_TEMPR4_2_net), .B(QX_TEMPR5_2_net), .S(BUFF_2_Y), 
        .Y(MX2_69_Y));
    BUFF BUFF_4 (.A(ADDRB_FF2_0_net), .Y(BUFF_4_Y));
    MX2 MX2_151 (.A(QX_TEMPR2_2_net), .B(QX_TEMPR3_2_net), .S(BUFF_2_Y)
        , .Y(MX2_151_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R6C0.mem") )  RAM_R6C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_6_net), .WEN(BLKA_EN_6_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R6C0_RD17), .RD16(RAM_R6C0_RD16), .RD15(
        RAM_R6C0_RD15), .RD14(RAM_R6C0_RD14), .RD13(RAM_R6C0_RD13), 
        .RD12(RAM_R6C0_RD12), .RD11(QX_TEMPR6_11_net), .RD10(
        QX_TEMPR6_10_net), .RD9(QX_TEMPR6_9_net), .RD8(QX_TEMPR6_8_net)
        , .RD7(QX_TEMPR6_7_net), .RD6(QX_TEMPR6_6_net), .RD5(
        QX_TEMPR6_5_net), .RD4(QX_TEMPR6_4_net), .RD3(QX_TEMPR6_3_net), 
        .RD2(QX_TEMPR6_2_net), .RD1(QX_TEMPR6_1_net), .RD0(
        QX_TEMPR6_0_net));
    MX2 MX2_RD_11_inst_inst_1 (.A(MX2_154_Y), .B(MX2_58_Y), .S(
        BUFF_9_Y), .Y(MX2_RD_11_inst));
    MX2 MX2_4 (.A(QX_TEMPR0_9_net), .B(QX_TEMPR1_9_net), .S(BUFF_1_Y), 
        .Y(MX2_4_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R3C0.mem") )  RAM_R3C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_3_net), .WEN(BLKA_EN_3_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R3C0_RD17), .RD16(RAM_R3C0_RD16), .RD15(
        RAM_R3C0_RD15), .RD14(RAM_R3C0_RD14), .RD13(RAM_R3C0_RD13), 
        .RD12(RAM_R3C0_RD12), .RD11(QX_TEMPR3_11_net), .RD10(
        QX_TEMPR3_10_net), .RD9(QX_TEMPR3_9_net), .RD8(QX_TEMPR3_8_net)
        , .RD7(QX_TEMPR3_7_net), .RD6(QX_TEMPR3_6_net), .RD5(
        QX_TEMPR3_5_net), .RD4(QX_TEMPR3_4_net), .RD3(QX_TEMPR3_3_net), 
        .RD2(QX_TEMPR3_2_net), .RD1(QX_TEMPR3_1_net), .RD0(
        QX_TEMPR3_0_net));
    NAND2 NAND2_ENABLE_ADDRB_2_inst (.A(AND2A_7_Y), .B(NOR2_3_Y), .Y(
        ENABLE_ADDRB_2_net));
    MX2 MX2_79 (.A(QX_TEMPR14_11_net), .B(QX_TEMPR15_11_net), .S(
        BUFF_7_Y), .Y(MX2_79_Y));
    MX2 MX2_43 (.A(QX_TEMPR10_2_net), .B(QX_TEMPR11_2_net), .S(
        BUFF_2_Y), .Y(MX2_43_Y));
    DFN1 BFF1_3_inst (.D(addr[11]), .CLK(n_rdclk), .Q(ADDRB_FF2_3_net));
    MX2 MX2_50 (.A(MX2_145_Y), .B(MX2_97_Y), .S(BUFF_10_Y), .Y(
        MX2_50_Y));
    BUFF BUFF_13 (.A(ADDRB_FF2_0_net), .Y(BUFF_13_Y));
    RAM512X18 #( .MEMORYFILE("RAM_R10C0.mem") )  RAM_R10C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_10_net), .WEN(BLKA_EN_10_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R10C0_RD17), .RD16(RAM_R10C0_RD16), .RD15(
        RAM_R10C0_RD15), .RD14(RAM_R10C0_RD14), .RD13(RAM_R10C0_RD13), 
        .RD12(RAM_R10C0_RD12), .RD11(QX_TEMPR10_11_net), .RD10(
        QX_TEMPR10_10_net), .RD9(QX_TEMPR10_9_net), .RD8(
        QX_TEMPR10_8_net), .RD7(QX_TEMPR10_7_net), .RD6(
        QX_TEMPR10_6_net), .RD5(QX_TEMPR10_5_net), .RD4(
        QX_TEMPR10_4_net), .RD3(QX_TEMPR10_3_net), .RD2(
        QX_TEMPR10_2_net), .RD1(QX_TEMPR10_1_net), .RD0(
        QX_TEMPR10_0_net));
    MX2 MX2_145 (.A(MX2_4_Y), .B(MX2_104_Y), .S(BUFF_18_Y), .Y(
        MX2_145_Y));
    MX2 MX2_103 (.A(MX2_59_Y), .B(MX2_120_Y), .S(BUFF_18_Y), .Y(
        MX2_103_Y));
    MX2 MX2_64 (.A(QX_TEMPR0_0_net), .B(QX_TEMPR1_0_net), .S(BUFF_11_Y)
        , .Y(MX2_64_Y));
    MX2 MX2_12 (.A(QX_TEMPR8_5_net), .B(QX_TEMPR9_5_net), .S(BUFF_12_Y)
        , .Y(MX2_12_Y));
    MX2 MX2_39 (.A(MX2_53_Y), .B(MX2_8_Y), .S(BUFF_16_Y), .Y(MX2_39_Y));
    NAND2 NAND2_ENABLE_ADDRB_0_inst (.A(NOR2_0_Y), .B(NOR2_3_Y), .Y(
        ENABLE_ADDRB_0_net));
    MX2 MX2_74 (.A(QX_TEMPR14_9_net), .B(QX_TEMPR15_9_net), .S(
        BUFF_6_Y), .Y(MX2_74_Y));
    MX2 MX2_167 (.A(QX_TEMPR2_10_net), .B(QX_TEMPR3_10_net), .S(
        BUFF_6_Y), .Y(MX2_167_Y));
    MX2 MX2_81 (.A(MX2_135_Y), .B(MX2_28_Y), .S(BUFF_10_Y), .Y(
        MX2_81_Y));
    MX2 MX2_101 (.A(QX_TEMPR8_7_net), .B(QX_TEMPR9_7_net), .S(BUFF_4_Y)
        , .Y(MX2_101_Y));
    OR2 ORB_GATE_11_inst (.A(ENABLE_ADDRB_11_net), .B(WEBP), .Y(
        BLKB_EN_11_net));
    MX2 MX2_122 (.A(MX2_73_Y), .B(MX2_21_Y), .S(BUFF_15_Y), .Y(
        MX2_122_Y));
    OR2 ORB_GATE_3_inst (.A(ENABLE_ADDRB_3_net), .B(WEBP), .Y(
        BLKB_EN_3_net));
    MX2 MX2_99 (.A(QX_TEMPR6_3_net), .B(QX_TEMPR7_3_net), .S(BUFF_13_Y)
        , .Y(MX2_99_Y));
    MX2 MX2_47 (.A(QX_TEMPR10_10_net), .B(QX_TEMPR11_10_net), .S(
        BUFF_6_Y), .Y(MX2_47_Y));
    NAND2 NAND2_ENABLE_ADDRA_9_inst (.A(AND2A_2_Y), .B(AND2A_1_Y), .Y(
        ENABLE_ADDRA_9_net));
    MX2 MX2_34 (.A(MX2_161_Y), .B(MX2_108_Y), .S(BUFF_15_Y), .Y(
        MX2_34_Y));
    MX2 MX2_18 (.A(QX_TEMPR12_10_net), .B(QX_TEMPR13_10_net), .S(
        BUFF_7_Y), .Y(MX2_18_Y));
    MX2 MX2_138 (.A(MX2_19_Y), .B(MX2_99_Y), .S(BUFF_16_Y), .Y(
        MX2_138_Y));
    NAND2 NAND2_ENABLE_ADDRB_9_inst (.A(AND2A_6_Y), .B(AND2A_5_Y), .Y(
        ENABLE_ADDRB_9_net));
    NAND2 NAND2_ENABLE_ADDRB_5_inst (.A(AND2A_6_Y), .B(AND2A_3_Y), .Y(
        ENABLE_ADDRB_5_net));
    RAM512X18 #( .MEMORYFILE("RAM_R7C0.mem") )  RAM_R7C0 (.RADDR8(
        RAM_GND), .RADDR7(addr[7]), .RADDR6(addr[6]), .RADDR5(addr[5]), 
        .RADDR4(addr[4]), .RADDR3(addr[3]), .RADDR2(addr[2]), .RADDR1(
        addr[1]), .RADDR0(addr[0]), .WADDR8(RAM_GND), .WADDR7(
        addr_0[7]), .WADDR6(addr_0[6]), .WADDR5(addr_0[5]), .WADDR4(
        addr_0[4]), .WADDR3(addr_0[3]), .WADDR2(addr_0[2]), .WADDR1(
        addr_0[1]), .WADDR0(addr_0[0]), .WD17(RAM_GND), .WD16(RAM_GND), 
        .WD15(RAM_GND), .WD14(RAM_GND), .WD13(RAM_GND), .WD12(RAM_GND), 
        .WD11(un1_n_s_change_0[11]), .WD10(un1_n_s_change_0[10]), .WD9(
        un1_n_s_change_0[9]), .WD8(un1_n_s_change_0[8]), .WD7(
        un1_n_s_change_0[7]), .WD6(un1_n_s_change_0[6]), .WD5(
        un1_n_s_change_0[5]), .WD4(un1_n_s_change_0[4]), .WD3(
        un1_n_s_change_0[3]), .WD2(un1_n_s_change_0[2]), .WD1(
        un1_n_s_change_0[1]), .WD0(un1_n_s_change_0[0]), .RW0(RAM_GND), 
        .RW1(RAM_VCC), .WW0(RAM_GND), .WW1(RAM_VCC), .PIPE(RAM_GND), 
        .REN(BLKB_EN_7_net), .WEN(BLKA_EN_7_net), .RCLK(n_rdclk), 
        .WCLK(s_clk_div4_0_clkout), .RESET(n_acq_change_0_n_rst_n_0), 
        .RD17(RAM_R7C0_RD17), .RD16(RAM_R7C0_RD16), .RD15(
        RAM_R7C0_RD15), .RD14(RAM_R7C0_RD14), .RD13(RAM_R7C0_RD13), 
        .RD12(RAM_R7C0_RD12), .RD11(QX_TEMPR7_11_net), .RD10(
        QX_TEMPR7_10_net), .RD9(QX_TEMPR7_9_net), .RD8(QX_TEMPR7_8_net)
        , .RD7(QX_TEMPR7_7_net), .RD6(QX_TEMPR7_6_net), .RD5(
        QX_TEMPR7_5_net), .RD4(QX_TEMPR7_4_net), .RD3(QX_TEMPR7_3_net), 
        .RD2(QX_TEMPR7_2_net), .RD1(QX_TEMPR7_1_net), .RD0(
        QX_TEMPR7_0_net));
    BUFF BUFF_11 (.A(ADDRB_FF2_0_net), .Y(BUFF_11_Y));
    MX2 MX2_137 (.A(QX_TEMPR8_4_net), .B(QX_TEMPR9_4_net), .S(
        BUFF_14_Y), .Y(MX2_137_Y));
    NAND2 NAND2_ENABLE_ADDRA_10_inst (.A(AND2A_4_Y), .B(AND2A_1_Y), .Y(
        ENABLE_ADDRA_10_net));
    MX2 MX2_94 (.A(MX2_129_Y), .B(MX2_17_Y), .S(BUFF_3_Y), .Y(MX2_94_Y)
        );
    MX2 MX2_16 (.A(MX2_3_Y), .B(MX2_167_Y), .S(BUFF_5_Y), .Y(MX2_16_Y));
    NAND2 NAND2_ENABLE_ADDRB_1_inst (.A(AND2A_6_Y), .B(NOR2_3_Y), .Y(
        ENABLE_ADDRB_1_net));
    MX2 MX2_85 (.A(QX_TEMPR14_3_net), .B(QX_TEMPR15_3_net), .S(
        BUFF_13_Y), .Y(MX2_85_Y));
    OR2 ORA_GATE_3_inst (.A(ENABLE_ADDRA_3_net), .B(WEAP), .Y(
        BLKA_EN_3_net));
    BUFF BUFF_18 (.A(ADDRB_FF2_1_net), .Y(BUFF_18_Y));
    OR2 ORB_GATE_0_inst (.A(ENABLE_ADDRB_0_net), .B(WEBP), .Y(
        BLKB_EN_0_net));
    MX2 MX2_126 (.A(QX_TEMPR6_10_net), .B(QX_TEMPR7_10_net), .S(
        BUFF_6_Y), .Y(MX2_126_Y));
    BUFF BUFF_1 (.A(ADDRB_FF2_0_net), .Y(BUFF_1_Y));
    MX2 MX2_162 (.A(MX2_22_Y), .B(MX2_111_Y), .S(BUFF_18_Y), .Y(
        MX2_162_Y));
    MX2 MX2_1 (.A(QX_TEMPR10_6_net), .B(QX_TEMPR11_6_net), .S(
        BUFF_12_Y), .Y(MX2_1_Y));
    MX2 MX2_13 (.A(QX_TEMPR8_8_net), .B(QX_TEMPR9_8_net), .S(BUFF_1_Y), 
        .Y(MX2_13_Y));
    MX2 MX2_144 (.A(QX_TEMPR10_5_net), .B(QX_TEMPR11_5_net), .S(
        BUFF_12_Y), .Y(MX2_144_Y));
    NAND2 NAND2_ENABLE_ADDRA_8_inst (.A(NOR2_2_Y), .B(AND2A_1_Y), .Y(
        ENABLE_ADDRA_8_net));
    MX2 MX2_140 (.A(MX2_14_Y), .B(MX2_147_Y), .S(BUFF_17_Y), .Y(
        MX2_140_Y));
    DFN1 BFF1_2_inst (.D(addr[10]), .CLK(n_rdclk), .Q(ADDRB_FF2_2_net));
    MX2 MX2_149 (.A(MX2_75_Y), .B(MX2_127_Y), .S(BUFF_16_Y), .Y(
        MX2_149_Y));
    
endmodule


module noise_addr_noise_addr_0_1(
       addr,
       top_code_0_RAM_Rd_rst,
       n_rdclk
    );
output [11:0] addr;
input  top_code_0_RAM_Rd_rst;
input  n_rdclk;

    wire \un1_noise_addr_1_i[0] , addr_n11, addr_c9, addr_n10, addr_n9, 
        addr_c8, addr_n8, addr_c6, addr_n7, addr_n6, addr_c4, addr_n5, 
        addr_n4, addr_c2, addr_n3, addr_n2, addr_n1, GND, VCC, GND_0, 
        VCC_0;
    
    DFN0C0 \addr[6]  (.D(addr_n6), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[6]));
    DFN0C0 \addr[11]  (.D(addr_n11), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[11]));
    XNOR2 \addr_RNO[7]  (.A(addr[7]), .B(addr_c6), .Y(addr_n7));
    AX1 \addr_RNO[6]  (.A(addr_c4), .B(addr[5]), .C(addr[6]), .Y(
        addr_n6));
    XNOR2 \addr_RNO[3]  (.A(addr[3]), .B(addr_c2), .Y(addr_n3));
    NOR3B \addr_RNIKU152[8]  (.A(addr[7]), .B(addr[8]), .C(addr_c6), 
        .Y(addr_c8));
    XOR2 \addr_RNO[1]  (.A(addr[1]), .B(addr[0]), .Y(addr_n1));
    VCC VCC_i (.Y(VCC));
    DFN0C0 \addr[3]  (.D(addr_n3), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[3]));
    DFN0C0 \addr[8]  (.D(addr_n8), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[8]));
    INV \addr_RNO[0]  (.A(addr[0]), .Y(\un1_noise_addr_1_i[0] ));
    DFN0C0 \addr[9]  (.D(addr_n9), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[9]));
    XOR2 \addr_RNO[9]  (.A(addr[9]), .B(addr_c8), .Y(addr_n9));
    OR3C \addr_RNIJK0N[2]  (.A(addr[0]), .B(addr[1]), .C(addr[2]), .Y(
        addr_c2));
    DFN0C0 \addr[0]  (.D(\un1_noise_addr_1_i[0] ), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[0]));
    OR3B \addr_RNI5RML1[6]  (.A(addr[5]), .B(addr[6]), .C(addr_c4), .Y(
        addr_c6));
    DFN0C0 \addr[4]  (.D(addr_n4), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[4]));
    DFN0C0 \addr[5]  (.D(addr_n5), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[5]));
    GND GND_i (.Y(GND));
    NOR2B \addr_RNIDGNC2[9]  (.A(addr[9]), .B(addr_c8), .Y(addr_c9));
    AX1C \addr_RNO[2]  (.A(addr[0]), .B(addr[1]), .C(addr[2]), .Y(
        addr_n2));
    OR3B \addr_RNIQNB61[4]  (.A(addr[3]), .B(addr[4]), .C(addr_c2), .Y(
        addr_c4));
    AX1C \addr_RNO[11]  (.A(addr_c9), .B(addr[10]), .C(addr[11]), .Y(
        addr_n11));
    DFN0C0 \addr[2]  (.D(addr_n2), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[2]));
    XOR2 \addr_RNO[10]  (.A(addr[10]), .B(addr_c9), .Y(addr_n10));
    XNOR2 \addr_RNO[5]  (.A(addr[5]), .B(addr_c4), .Y(addr_n5));
    DFN0C0 \addr[10]  (.D(addr_n10), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[10]));
    DFN0C0 \addr[7]  (.D(addr_n7), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[7]));
    AX1 \addr_RNO[4]  (.A(addr_c2), .B(addr[3]), .C(addr[4]), .Y(
        addr_n4));
    DFN0C0 \addr[1]  (.D(addr_n1), .CLK(n_rdclk), .CLR(
        top_code_0_RAM_Rd_rst), .Q(addr[1]));
    AX1 \addr_RNO[8]  (.A(addr_c6), .B(addr[7]), .C(addr[8]), .Y(
        addr_n8));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module noise_acq(
       un1_n_s_change_0,
       n_acqnum,
       n_divnum,
       top_code_0_RAM_Rd_rst,
       MX2_RD_0_inst,
       MX2_RD_2_inst,
       noise_acq_GND,
       noise_acq_VCC,
       MX2_RD_4_inst,
       MX2_RD_5_inst,
       MX2_RD_7_inst,
       MX2_RD_6_inst,
       MX2_RD_11_inst,
       MX2_RD_1_inst,
       MX2_RD_9_inst,
       MX2_RD_3_inst,
       MX2_RD_10_inst,
       MX2_RD_8_inst,
       n_acq_change_0_n_acq_start,
       top_code_0_n_load,
       s_clk_div4_0_clkout,
       n_acq_change_0_n_rst_n,
       top_code_0_n_rd_en,
       n_acq_change_0_n_rst_n_0,
       XRD_c,
       GLA
    );
input  [11:0] un1_n_s_change_0;
input  [11:0] n_acqnum;
input  [9:0] n_divnum;
input  top_code_0_RAM_Rd_rst;
output MX2_RD_0_inst;
output MX2_RD_2_inst;
input  noise_acq_GND;
input  noise_acq_VCC;
output MX2_RD_4_inst;
output MX2_RD_5_inst;
output MX2_RD_7_inst;
output MX2_RD_6_inst;
output MX2_RD_11_inst;
output MX2_RD_1_inst;
output MX2_RD_9_inst;
output MX2_RD_3_inst;
output MX2_RD_10_inst;
output MX2_RD_8_inst;
input  n_acq_change_0_n_acq_start;
input  top_code_0_n_load;
output s_clk_div4_0_clkout;
input  n_acq_change_0_n_rst_n;
input  top_code_0_n_rd_en;
input  n_acq_change_0_n_rst_n_0;
input  XRD_c;
input  GLA;

    wire n_rdclk, \addr_0[0] , \addr_0[1] , \addr_0[2] , \addr_0[3] , 
        \addr_0[4] , \addr_0[5] , \addr_0[6] , \addr_0[7] , 
        \addr_0[8] , \addr_0[9] , \addr_0[10] , \addr_0[11] , 
        noiseclkctrl_0_en, \addr[0] , \addr[1] , \addr[2] , \addr[3] , 
        \addr[4] , \addr[5] , \addr[6] , \addr[7] , \addr[8] , 
        \addr[9] , \addr[10] , \addr[11] , GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    n_rdclk_syn n_rdclk_syn_0 (.n_rdclk(n_rdclk), .GLA(GLA), .XRD_c(
        XRD_c), .n_acq_change_0_n_rst_n_0(n_acq_change_0_n_rst_n_0), 
        .top_code_0_n_rd_en(top_code_0_n_rd_en));
    noise_addr_noise_addr_0 noise_addr_0 (.addr_0({\addr_0[11] , 
        \addr_0[10] , \addr_0[9] , \addr_0[8] , \addr_0[7] , 
        \addr_0[6] , \addr_0[5] , \addr_0[4] , \addr_0[3] , 
        \addr_0[2] , \addr_0[1] , \addr_0[0] }), 
        .n_acq_change_0_n_rst_n(n_acq_change_0_n_rst_n), 
        .n_acq_change_0_n_rst_n_0(n_acq_change_0_n_rst_n_0), 
        .s_clk_div4_0_clkout(s_clk_div4_0_clkout));
    GND GND_i_0 (.Y(GND_0));
    noiseclk noiseclk_0 (.n_divnum({n_divnum[9], n_divnum[8], 
        n_divnum[7], n_divnum[6], n_divnum[5], n_divnum[4], 
        n_divnum[3], n_divnum[2], n_divnum[1], n_divnum[0]}), 
        .top_code_0_n_load(top_code_0_n_load), .GLA(GLA), 
        .s_clk_div4_0_clkout(s_clk_div4_0_clkout), .noiseclkctrl_0_en(
        noiseclkctrl_0_en), .n_acq_change_0_n_acq_start(
        n_acq_change_0_n_acq_start), .n_acq_change_0_n_rst_n_0(
        n_acq_change_0_n_rst_n_0));
    noiseclkctrl noiseclkctrl_0 (.n_acqnum({n_acqnum[11], n_acqnum[10], 
        n_acqnum[9], n_acqnum[8], n_acqnum[7], n_acqnum[6], 
        n_acqnum[5], n_acqnum[4], n_acqnum[3], n_acqnum[2], 
        n_acqnum[1], n_acqnum[0]}), .top_code_0_n_load(
        top_code_0_n_load), .GLA(GLA), .n_acq_change_0_n_rst_n(
        n_acq_change_0_n_rst_n), .s_clk_div4_0_clkout(
        s_clk_div4_0_clkout), .noiseclkctrl_0_en(noiseclkctrl_0_en));
    VCC VCC_i (.Y(VCC));
    RAM RAM_0 (.un1_n_s_change_0({un1_n_s_change_0[11], 
        un1_n_s_change_0[10], un1_n_s_change_0[9], un1_n_s_change_0[8], 
        un1_n_s_change_0[7], un1_n_s_change_0[6], un1_n_s_change_0[5], 
        un1_n_s_change_0[4], un1_n_s_change_0[3], un1_n_s_change_0[2], 
        un1_n_s_change_0[1], un1_n_s_change_0[0]}), .addr_0({
        \addr_0[11] , \addr_0[10] , \addr_0[9] , \addr_0[8] , 
        \addr_0[7] , \addr_0[6] , \addr_0[5] , \addr_0[4] , 
        \addr_0[3] , \addr_0[2] , \addr_0[1] , \addr_0[0] }), .addr({
        \addr[11] , \addr[10] , \addr[9] , \addr[8] , \addr[7] , 
        \addr[6] , \addr[5] , \addr[4] , \addr[3] , \addr[2] , 
        \addr[1] , \addr[0] }), .MX2_RD_8_inst(MX2_RD_8_inst), 
        .MX2_RD_10_inst(MX2_RD_10_inst), .MX2_RD_3_inst(MX2_RD_3_inst), 
        .MX2_RD_9_inst(MX2_RD_9_inst), .MX2_RD_1_inst(MX2_RD_1_inst), 
        .top_code_0_n_rd_en(top_code_0_n_rd_en), .MX2_RD_11_inst(
        MX2_RD_11_inst), .MX2_RD_6_inst(MX2_RD_6_inst), .MX2_RD_7_inst(
        MX2_RD_7_inst), .n_acq_change_0_n_acq_start(
        n_acq_change_0_n_acq_start), .MX2_RD_5_inst(MX2_RD_5_inst), 
        .MX2_RD_4_inst(MX2_RD_4_inst), .s_clk_div4_0_clkout(
        s_clk_div4_0_clkout), .RAM_VCC(noise_acq_VCC), 
        .n_acq_change_0_n_rst_n_0(n_acq_change_0_n_rst_n_0), .n_rdclk(
        n_rdclk), .RAM_GND(noise_acq_GND), .MX2_RD_2_inst(
        MX2_RD_2_inst), .MX2_RD_0_inst(MX2_RD_0_inst));
    noise_addr_noise_addr_0_1 noise_addr_1 (.addr({\addr[11] , 
        \addr[10] , \addr[9] , \addr[8] , \addr[7] , \addr[6] , 
        \addr[5] , \addr[4] , \addr[3] , \addr[2] , \addr[1] , 
        \addr[0] }), .top_code_0_RAM_Rd_rst(top_code_0_RAM_Rd_rst), 
        .n_rdclk(n_rdclk));
    GND GND_i (.Y(GND));
    
endmodule


module Signal_Noise_Acq(
       dataout_0,
       n_divnum,
       n_acqnum,
       s_addchoice,
       s_acqnum,
       s_periodnum,
       s_stripnum,
       ADC_c,
       Signal_Noise_Acq_0_acq_clk,
       XRD_c,
       n_acq_change_0_n_rst_n_0,
       top_code_0_n_rd_en,
       n_acq_change_0_n_rst_n,
       top_code_0_n_load,
       n_acq_change_0_n_acq_start,
       Signal_Noise_Acq_VCC,
       Signal_Noise_Acq_GND,
       top_code_0_RAM_Rd_rst,
       s_acq_change_0_s_rst,
       ddsclkout_c,
       scan_scale_sw_0_s_start,
       s_acq_change_0_s_load_0,
       s_acq_change_0_s_load,
       GLA,
       top_code_0_n_s_ctrl,
       top_code_0_n_s_ctrl_1,
       top_code_0_n_s_ctrl_0
    );
output [15:0] dataout_0;
input  [9:0] n_divnum;
input  [11:0] n_acqnum;
input  [4:0] s_addchoice;
input  [15:0] s_acqnum;
input  [3:0] s_periodnum;
input  [11:0] s_stripnum;
input  [11:0] ADC_c;
output Signal_Noise_Acq_0_acq_clk;
input  XRD_c;
input  n_acq_change_0_n_rst_n_0;
input  top_code_0_n_rd_en;
input  n_acq_change_0_n_rst_n;
input  top_code_0_n_load;
input  n_acq_change_0_n_acq_start;
input  Signal_Noise_Acq_VCC;
input  Signal_Noise_Acq_GND;
input  top_code_0_RAM_Rd_rst;
input  s_acq_change_0_s_rst;
input  ddsclkout_c;
input  scan_scale_sw_0_s_start;
input  s_acq_change_0_s_load_0;
input  s_acq_change_0_s_load;
input  GLA;
input  top_code_0_n_s_ctrl;
input  top_code_0_n_s_ctrl_1;
input  top_code_0_n_s_ctrl_0;

    wire \un1_n_s_change_0_1[11]_net_1 , 
        \un1_n_s_change_0_1[10]_net_1 , \un1_n_s_change_0[11]_net_1 , 
        \un1_n_s_change_0[10]_net_1 , \un1_n_s_change_0_1[6]_net_1 , 
        \un1_n_s_change_0_1[4]_net_1 , \un1_n_s_change_0[6]_net_1 , 
        \un1_n_s_change_0[4]_net_1 , \un1_n_s_change_0_1[9]_net_1 , 
        \un1_n_s_change_0_1[5]_net_1 , \un1_n_s_change_0_1[3]_net_1 , 
        \un1_n_s_change_0[9]_net_1 , \un1_n_s_change_0[5]_net_1 , 
        \un1_n_s_change_0[3]_net_1 , \un1_n_s_change_0[7]_net_1 , 
        \un1_n_s_change_0_1[7]_net_1 , \un1_n_s_change_0[8]_net_1 , 
        \un1_n_s_change_0_1[8]_net_1 , \un1_n_s_change_0[0]_net_1 , 
        \un1_n_s_change_0_1[0]_net_1 , \un1_n_s_change_0[1]_net_1 , 
        \un1_n_s_change_0_1[1]_net_1 , \un1_n_s_change_0_1[2]_net_1 , 
        \un1_n_s_change_0[2]_net_1 , \un1_add_reg_4_i[13] , 
        \un1_add_reg_4_i[15] , \addresult_0[13] , \addresult_0[15] , 
        \addresult_RNIJE5C[14] , \addresult[12] , \addresult[13] , 
        \addresult[14] , \addresult[15] , \un1_signal_acq_0[0] , 
        \un1_signal_acq_0[1] , \un1_signal_acq_0[2] , 
        \un1_signal_acq_0[3] , \addresult_4[13] , \addresult_4[15] , 
        \addresult_RNI8MQ7[14] , \addresult_5[13] , \addresult_5[15] , 
        \addresult_RNI7DQA[14] , \addresult_RNI5DQA[12] , N_104, N_88, 
        N_86, N_27_i_0, N_22_i_0, N_18_i_0, N_16_i_0, N_14_i_0, 
        N_12_i_0, N_20_i_0, N_25_i_0, N_92, N_108, N_99, N_115, N_107, 
        N_91, N_97, N_113, N_105, N_89, N_87, N_95, N_111, 
        signal_acq_0_Signal_acq_clk, N_33, N_256, N_255, N_253, N_251, 
        N_39, MX2_RD_0_inst, MX2_RD_2_inst, MX2_RD_4_inst, 
        MX2_RD_5_inst, MX2_RD_7_inst, MX2_RD_6_inst, MX2_RD_11_inst, 
        MX2_RD_1_inst, MX2_RD_9_inst, MX2_RD_3_inst, MX2_RD_10_inst, 
        MX2_RD_8_inst, s_clk_div4_0_clkout, GND, VCC, GND_0, VCC_0;
    
    OR2A \un1_n_s_change_0_1[4]  (.A(ADC_c[4]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[4]_net_1 ));
    NOR2B \un1_n_s_change_0[8]  (.A(top_code_0_n_s_ctrl), .B(ADC_c[8]), 
        .Y(\un1_n_s_change_0[8]_net_1 ));
    OR2A \un1_n_s_change_0_1[6]  (.A(ADC_c[6]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[6]_net_1 ));
    OR2A \un1_n_s_change_0_1[1]  (.A(ADC_c[1]), .B(top_code_0_n_s_ctrl)
        , .Y(\un1_n_s_change_0_1[1]_net_1 ));
    NOR2A \un1_n_s_change_0_1[5]  (.A(ADC_c[5]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[5]_net_1 ));
    NOR2B \un1_n_s_change_0[6]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[6]), .Y(\un1_n_s_change_0[6]_net_1 ));
    OR2A \un1_n_s_change_0_1[3]  (.A(ADC_c[3]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[3]_net_1 ));
    OR2A \un1_n_s_change_0_1[10]  (.A(ADC_c[10]), .B(
        top_code_0_n_s_ctrl_0), .Y(\un1_n_s_change_0_1[10]_net_1 ));
    OR2A \un1_n_s_change_0_1[2]  (.A(ADC_c[2]), .B(top_code_0_n_s_ctrl)
        , .Y(\un1_n_s_change_0_1[2]_net_1 ));
    NOR2B \un1_n_s_change_0[0]  (.A(top_code_0_n_s_ctrl), .B(ADC_c[0]), 
        .Y(\un1_n_s_change_0[0]_net_1 ));
    GND GND_i_0 (.Y(GND_0));
    OR2A \un1_n_s_change_0_1[9]  (.A(ADC_c[9]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[9]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR2B \un1_n_s_change_0[3]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[3]), .Y(\un1_n_s_change_0[3]_net_1 ));
    NOR2B \un1_n_s_change_0[1]  (.A(top_code_0_n_s_ctrl), .B(ADC_c[1]), 
        .Y(\un1_n_s_change_0[1]_net_1 ));
    OR2A \un1_n_s_change_0_1[11]  (.A(ADC_c[11]), .B(
        top_code_0_n_s_ctrl_0), .Y(\un1_n_s_change_0_1[11]_net_1 ));
    NOR2B \un1_n_s_change_0[5]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[5]), .Y(\un1_n_s_change_0[5]_net_1 ));
    OR2A \un1_n_s_change_0_1[0]  (.A(ADC_c[0]), .B(top_code_0_n_s_ctrl)
        , .Y(\un1_n_s_change_0_1[0]_net_1 ));
    GND GND_i (.Y(GND));
    NOR2B \un1_n_s_change_0[11]  (.A(top_code_0_n_s_ctrl_0), .B(
        ADC_c[11]), .Y(\un1_n_s_change_0[11]_net_1 ));
    NOR2B \un1_n_s_change_0[10]  (.A(top_code_0_n_s_ctrl_0), .B(
        ADC_c[10]), .Y(\un1_n_s_change_0[10]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2B \un1_n_s_change_0[9]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[9]), .Y(\un1_n_s_change_0[9]_net_1 ));
    signal_acq signal_acq_0 (.un1_add_reg_4_i_0(\un1_add_reg_4_i[13] ), 
        .un1_add_reg_4_i_2(\un1_add_reg_4_i[15] ), .ADC_c({ADC_c[2], 
        ADC_c[1], ADC_c[0]}), .addresult_0_0(\addresult_0[13] ), 
        .addresult_0_2(\addresult_0[15] ), .addresult_RNIJE5C({
        \addresult_RNIJE5C[14] }), .addresult({\addresult[15] , 
        \addresult[14] , \addresult[13] , \addresult[12] }), 
        .un1_signal_acq_0({\un1_signal_acq_0[3] , 
        \un1_signal_acq_0[2] , \un1_signal_acq_0[1] , 
        \un1_signal_acq_0[0] }), .addresult_4_0(\addresult_4[13] ), 
        .addresult_4_2(\addresult_4[15] ), .addresult_RNI8MQ7({
        \addresult_RNI8MQ7[14] }), .s_stripnum({s_stripnum[11], 
        s_stripnum[10], s_stripnum[9], s_stripnum[8], s_stripnum[7], 
        s_stripnum[6], s_stripnum[5], s_stripnum[4], s_stripnum[3], 
        s_stripnum[2], s_stripnum[1], s_stripnum[0]}), .s_periodnum({
        s_periodnum[3], s_periodnum[2], s_periodnum[1], s_periodnum[0]})
        , .s_acqnum({s_acqnum[15], s_acqnum[14], s_acqnum[13], 
        s_acqnum[12], s_acqnum[11], s_acqnum[10], s_acqnum[9], 
        s_acqnum[8], s_acqnum[7], s_acqnum[6], s_acqnum[5], 
        s_acqnum[4], s_acqnum[3], s_acqnum[2], s_acqnum[1], 
        s_acqnum[0]}), .un1_n_s_change_0_1({
        \un1_n_s_change_0_1[11]_net_1 , \un1_n_s_change_0_1[10]_net_1 , 
        \un1_n_s_change_0_1[9]_net_1 , \un1_n_s_change_0_1[8]_net_1 , 
        \un1_n_s_change_0_1[7]_net_1 , \un1_n_s_change_0_1[6]_net_1 , 
        \un1_n_s_change_0_1[5]_net_1 , \un1_n_s_change_0_1[4]_net_1 , 
        \un1_n_s_change_0_1[3]_net_1 , \un1_n_s_change_0_1[2]_net_1 , 
        \un1_n_s_change_0_1[1]_net_1 , \un1_n_s_change_0_1[0]_net_1 }), 
        .addresult_5_0(\addresult_5[13] ), .addresult_5_2(
        \addresult_5[15] ), .addresult_RNI7DQA({
        \addresult_RNI7DQA[14] }), .addresult_RNI5DQA({
        \addresult_RNI5DQA[12] }), .s_addchoice({s_addchoice[4], 
        s_addchoice[3], s_addchoice[2], s_addchoice[1], s_addchoice[0]})
        , .top_code_0_n_s_ctrl_0(top_code_0_n_s_ctrl_0), .N_104(N_104), 
        .N_88(N_88), .N_86(N_86), .N_27_i_0(N_27_i_0), .N_22_i_0(
        N_22_i_0), .N_18_i_0(N_18_i_0), .N_16_i_0(N_16_i_0), .N_14_i_0(
        N_14_i_0), .N_12_i_0(N_12_i_0), .N_20_i_0(N_20_i_0), .N_25_i_0(
        N_25_i_0), .N_92(N_92), .N_108(N_108), .N_99(N_99), .N_115(
        N_115), .N_107(N_107), .N_91(N_91), .N_97(N_97), .N_113(N_113), 
        .N_105(N_105), .N_89(N_89), .N_87(N_87), .N_95(N_95), .N_111(
        N_111), .signal_acq_0_Signal_acq_clk(
        signal_acq_0_Signal_acq_clk), .GLA(GLA), 
        .s_acq_change_0_s_load(s_acq_change_0_s_load), 
        .s_acq_change_0_s_load_0(s_acq_change_0_s_load_0), 
        .scan_scale_sw_0_s_start(scan_scale_sw_0_s_start), 
        .ddsclkout_c(ddsclkout_c), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .N_33(N_33), .N_256(N_256), .N_255(
        N_255), .N_253(N_253), .N_251(N_251), .N_39(N_39));
    NOR2B \un1_n_s_change_0[2]  (.A(top_code_0_n_s_ctrl), .B(ADC_c[2]), 
        .Y(\un1_n_s_change_0[2]_net_1 ));
    OR2A \un1_n_s_change_0_1[8]  (.A(ADC_c[8]), .B(top_code_0_n_s_ctrl)
        , .Y(\un1_n_s_change_0_1[8]_net_1 ));
    NOR2B \un1_n_s_change_0[7]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[7]), .Y(\un1_n_s_change_0[7]_net_1 ));
    NOR2B \un1_n_s_change_0[4]  (.A(top_code_0_n_s_ctrl_1), .B(
        ADC_c[4]), .Y(\un1_n_s_change_0[4]_net_1 ));
    OR2A \un1_n_s_change_0_1[7]  (.A(ADC_c[7]), .B(
        top_code_0_n_s_ctrl_1), .Y(\un1_n_s_change_0_1[7]_net_1 ));
    n_s_change n_s_change_0 (.un1_signal_acq_0({\un1_signal_acq_0[3] , 
        \un1_signal_acq_0[2] , \un1_signal_acq_0[1] , 
        \un1_signal_acq_0[0] }), .dataout_0_2(dataout_0[2]), 
        .dataout_0_3(dataout_0[3]), .dataout_0_1(dataout_0[1]), 
        .dataout_0_5(dataout_0[5]), .dataout_0_11(dataout_0[11]), 
        .dataout_0_7(dataout_0[7]), .dataout_0_8(dataout_0[8]), 
        .dataout_0_6(dataout_0[6]), .dataout_0_0_d0(dataout_0[0]), 
        .dataout_0_10(dataout_0[10]), .dataout_0_9(dataout_0[9]), 
        .dataout_0_4(dataout_0[4]), .dataout_0_0({dataout_0[15], 
        dataout_0[14], dataout_0[13], dataout_0[12]}), 
        .addresult_RNI5DQA({\addresult_RNI5DQA[12] }), 
        .addresult_RNIJE5C({\addresult_RNIJE5C[14] }), 
        .addresult_RNI8MQ7({\addresult_RNI8MQ7[14] }), 
        .addresult_RNI7DQA({\addresult_RNI7DQA[14] }), .addresult({
        \addresult[15] , \addresult[14] , \addresult[13] , 
        \addresult[12] }), .addresult_0_0(\addresult_0[13] ), 
        .addresult_0_2(\addresult_0[15] ), .un1_add_reg_4_i_0(
        \un1_add_reg_4_i[13] ), .un1_add_reg_4_i_2(
        \un1_add_reg_4_i[15] ), .addresult_5_0(\addresult_5[13] ), 
        .addresult_5_2(\addresult_5[15] ), .addresult_4_0(
        \addresult_4[13] ), .addresult_4_2(\addresult_4[15] ), 
        .MX2_RD_2_inst(MX2_RD_2_inst), .MX2_RD_3_inst(MX2_RD_3_inst), 
        .MX2_RD_1_inst(MX2_RD_1_inst), .MX2_RD_5_inst(MX2_RD_5_inst), 
        .N_25_i_0(N_25_i_0), .top_code_0_n_s_ctrl(top_code_0_n_s_ctrl), 
        .MX2_RD_11_inst(MX2_RD_11_inst), .N_20_i_0(N_20_i_0), 
        .MX2_RD_7_inst(MX2_RD_7_inst), .N_12_i_0(N_12_i_0), 
        .s_clk_div4_0_clkout(s_clk_div4_0_clkout), 
        .signal_acq_0_Signal_acq_clk(signal_acq_0_Signal_acq_clk), 
        .Signal_Noise_Acq_0_acq_clk(Signal_Noise_Acq_0_acq_clk), 
        .top_code_0_n_s_ctrl_1(top_code_0_n_s_ctrl_1), .MX2_RD_8_inst(
        MX2_RD_8_inst), .N_14_i_0(N_14_i_0), .MX2_RD_6_inst(
        MX2_RD_6_inst), .N_27_i_0(N_27_i_0), .MX2_RD_0_inst(
        MX2_RD_0_inst), .MX2_RD_10_inst(MX2_RD_10_inst), .N_18_i_0(
        N_18_i_0), .MX2_RD_9_inst(MX2_RD_9_inst), .N_16_i_0(N_16_i_0), 
        .MX2_RD_4_inst(MX2_RD_4_inst), .N_22_i_0(N_22_i_0), .N_89(N_89)
        , .N_88(N_88), .N_92(N_92), .N_86(N_86), .N_87(N_87), .N_91(
        N_91), .N_95(N_95), .N_97(N_97), .N_99(N_99), .N_105(N_105), 
        .N_104(N_104), .N_108(N_108), .N_107(N_107), .N_33(N_33), 
        .N_256(N_256), .N_111(N_111), .N_255(N_255), .N_113(N_113), 
        .N_253(N_253), .N_115(N_115), .N_251(N_251), 
        .top_code_0_n_s_ctrl_0(top_code_0_n_s_ctrl_0), .N_39(N_39));
    noise_acq noise_acq_0 (.un1_n_s_change_0({
        \un1_n_s_change_0[11]_net_1 , \un1_n_s_change_0[10]_net_1 , 
        \un1_n_s_change_0[9]_net_1 , \un1_n_s_change_0[8]_net_1 , 
        \un1_n_s_change_0[7]_net_1 , \un1_n_s_change_0[6]_net_1 , 
        \un1_n_s_change_0[5]_net_1 , \un1_n_s_change_0[4]_net_1 , 
        \un1_n_s_change_0[3]_net_1 , \un1_n_s_change_0[2]_net_1 , 
        \un1_n_s_change_0[1]_net_1 , \un1_n_s_change_0[0]_net_1 }), 
        .n_acqnum({n_acqnum[11], n_acqnum[10], n_acqnum[9], 
        n_acqnum[8], n_acqnum[7], n_acqnum[6], n_acqnum[5], 
        n_acqnum[4], n_acqnum[3], n_acqnum[2], n_acqnum[1], 
        n_acqnum[0]}), .n_divnum({n_divnum[9], n_divnum[8], 
        n_divnum[7], n_divnum[6], n_divnum[5], n_divnum[4], 
        n_divnum[3], n_divnum[2], n_divnum[1], n_divnum[0]}), 
        .top_code_0_RAM_Rd_rst(top_code_0_RAM_Rd_rst), .MX2_RD_0_inst(
        MX2_RD_0_inst), .MX2_RD_2_inst(MX2_RD_2_inst), .noise_acq_GND(
        Signal_Noise_Acq_GND), .noise_acq_VCC(Signal_Noise_Acq_VCC), 
        .MX2_RD_4_inst(MX2_RD_4_inst), .MX2_RD_5_inst(MX2_RD_5_inst), 
        .MX2_RD_7_inst(MX2_RD_7_inst), .MX2_RD_6_inst(MX2_RD_6_inst), 
        .MX2_RD_11_inst(MX2_RD_11_inst), .MX2_RD_1_inst(MX2_RD_1_inst), 
        .MX2_RD_9_inst(MX2_RD_9_inst), .MX2_RD_3_inst(MX2_RD_3_inst), 
        .MX2_RD_10_inst(MX2_RD_10_inst), .MX2_RD_8_inst(MX2_RD_8_inst), 
        .n_acq_change_0_n_acq_start(n_acq_change_0_n_acq_start), 
        .top_code_0_n_load(top_code_0_n_load), .s_clk_div4_0_clkout(
        s_clk_div4_0_clkout), .n_acq_change_0_n_rst_n(
        n_acq_change_0_n_rst_n), .top_code_0_n_rd_en(
        top_code_0_n_rd_en), .n_acq_change_0_n_rst_n_0(
        n_acq_change_0_n_rst_n_0), .XRD_c(XRD_c), .GLA(GLA));
    
endmodule


module bri_dump_sw(
       bri_dump_sw_0_dump_start,
       bri_dump_sw_0_dumpoff_ctr,
       bri_dump_sw_0_off_test,
       bri_dump_sw_0_phase_ctr,
       pulse_start_c,
       bri_dump_sw_0_reset_out,
       bri_dump_sw_0_tetw_pluse,
       net_45,
       top_code_0_pluse_rst,
       scalestate_0_tetw_pluse,
       scalestate_0_pluse_start,
       scalestate_0_pn_out,
       top_code_0_pn_change,
       scalestate_0_off_test,
       plusestate_0_off_test,
       scalestate_0_dumpoff_ctr,
       plusestate_0_tetw_pluse,
       top_code_0_pluse_scale,
       scalestate_0_dump_start,
       plusestate_0_soft_d,
       net_27,
       GLA,
       bri_dump_sw_0_reset_out_0
    );
output bri_dump_sw_0_dump_start;
output bri_dump_sw_0_dumpoff_ctr;
output bri_dump_sw_0_off_test;
output bri_dump_sw_0_phase_ctr;
output pulse_start_c;
output bri_dump_sw_0_reset_out;
output bri_dump_sw_0_tetw_pluse;
input  net_45;
input  top_code_0_pluse_rst;
input  scalestate_0_tetw_pluse;
input  scalestate_0_pluse_start;
input  scalestate_0_pn_out;
input  top_code_0_pn_change;
input  scalestate_0_off_test;
input  plusestate_0_off_test;
input  scalestate_0_dumpoff_ctr;
input  plusestate_0_tetw_pluse;
input  top_code_0_pluse_scale;
input  scalestate_0_dump_start;
input  plusestate_0_soft_d;
input  net_27;
input  GLA;
output bri_dump_sw_0_reset_out_0;

    wire reset_out_0_net_1, tetw_pluse_RNO_net_1, tetw_pluse_5, 
        reset_out_5_net_1, pluse_start_RNO_0_net_1, pluse_start_5, 
        phase_ctr_RNO_net_1, phase_ctr_5, off_test_RNO_net_1, 
        off_test_5, dumpoff_ctr_RNO_0_net_1, dumpoff_ctr_5, 
        dump_start_RNO_0_net_1, dump_start_5, GND, VCC, GND_0, VCC_0;
    
    NOR2A phase_ctr_RNO (.A(net_27), .B(phase_ctr_5), .Y(
        phase_ctr_RNO_net_1));
    NOR2A tetw_pluse_RNO (.A(net_27), .B(tetw_pluse_5), .Y(
        tetw_pluse_RNO_net_1));
    DFN1 dump_start (.D(dump_start_RNO_0_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_dump_start));
    GND GND_i_0 (.Y(GND_0));
    MX2C reset_out_5 (.A(top_code_0_pluse_rst), .B(net_45), .S(
        top_code_0_pluse_scale), .Y(reset_out_5_net_1));
    MX2C pluse_start_RNO_0 (.A(plusestate_0_off_test), .B(
        scalestate_0_pluse_start), .S(top_code_0_pluse_scale), .Y(
        pluse_start_5));
    DFN1 off_test (.D(off_test_RNO_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_off_test));
    VCC VCC_i (.Y(VCC));
    MX2C off_test_RNO_0 (.A(plusestate_0_off_test), .B(
        scalestate_0_off_test), .S(top_code_0_pluse_scale), .Y(
        off_test_5));
    NOR2A dumpoff_ctr_RNO (.A(net_27), .B(dumpoff_ctr_5), .Y(
        dumpoff_ctr_RNO_0_net_1));
    MX2C phase_ctr_RNO_0 (.A(top_code_0_pn_change), .B(
        scalestate_0_pn_out), .S(top_code_0_pluse_scale), .Y(
        phase_ctr_5));
    DFN1 phase_ctr (.D(phase_ctr_RNO_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_phase_ctr));
    NOR2A off_test_RNO (.A(net_27), .B(off_test_5), .Y(
        off_test_RNO_net_1));
    MX2C tetw_pluse_RNO_0 (.A(plusestate_0_tetw_pluse), .B(
        scalestate_0_tetw_pluse), .S(top_code_0_pluse_scale), .Y(
        tetw_pluse_5));
    DFN1 reset_out_0_0 (.D(reset_out_0_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_reset_out_0));
    GND GND_i (.Y(GND));
    MX2C dump_start_RNO_0 (.A(plusestate_0_soft_d), .B(
        scalestate_0_dump_start), .S(top_code_0_pluse_scale), .Y(
        dump_start_5));
    DFN1 tetw_pluse (.D(tetw_pluse_RNO_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_tetw_pluse));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 dumpoff_ctr (.D(dumpoff_ctr_RNO_0_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_dumpoff_ctr));
    MX2C dumpoff_ctr_RNO_0 (.A(plusestate_0_tetw_pluse), .B(
        scalestate_0_dumpoff_ctr), .S(top_code_0_pluse_scale), .Y(
        dumpoff_ctr_5));
    DFN1 pluse_start (.D(pluse_start_RNO_0_net_1), .CLK(GLA), .Q(
        pulse_start_c));
    NOR2A dump_start_RNO (.A(net_27), .B(dump_start_5), .Y(
        dump_start_RNO_0_net_1));
    NOR2A pluse_start_RNO (.A(net_27), .B(pluse_start_5), .Y(
        pluse_start_RNO_0_net_1));
    NOR2A reset_out_0 (.A(net_27), .B(reset_out_5_net_1), .Y(
        reset_out_0_net_1));
    DFN1 reset_out (.D(reset_out_0_net_1), .CLK(GLA), .Q(
        bri_dump_sw_0_reset_out));
    
endmodule


module dump_sustain_timer(
       dump_sustain_timer_0_start,
       clk_5K,
       AND2_1_Y,
       scalestate_0_dump_sustain_ctrl
    );
output dump_sustain_timer_0_start;
input  clk_5K;
input  AND2_1_Y;
input  scalestate_0_dump_sustain_ctrl;

    wire N_6, \count[0]_net_1 , \count[1]_net_1 , N_11, 
        start_RNO_net_1, \count[2]_net_1 , N_9, count_n0, N_8, GND, 
        VCC, GND_0, VCC_0;
    
    DFN1 \count[0]  (.D(count_n0), .CLK(clk_5K), .Q(\count[0]_net_1 ));
    DFN1 start (.D(start_RNO_net_1), .CLK(clk_5K), .Q(
        dump_sustain_timer_0_start));
    XA1B \count_RNO[2]  (.A(N_9), .B(\count[2]_net_1 ), .C(N_11), .Y(
        N_8));
    DFN1 \count[2]  (.D(N_8), .CLK(clk_5K), .Q(\count[2]_net_1 ));
    NOR2 \count_RNO[0]  (.A(\count[0]_net_1 ), .B(N_11), .Y(count_n0));
    DFN1 \count[1]  (.D(N_6), .CLK(clk_5K), .Q(\count[1]_net_1 ));
    XA1B \count_RNO[1]  (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(N_11), .Y(N_6));
    VCC VCC_i_0 (.Y(VCC_0));
    VCC VCC_i (.Y(VCC));
    NOR3C start_RNO (.A(\count[2]_net_1 ), .B(
        scalestate_0_dump_sustain_ctrl), .C(N_9), .Y(start_RNO_net_1));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    NOR2B \count_RNI9I5E[1]  (.A(\count[1]_net_1 ), .B(
        \count[0]_net_1 ), .Y(N_9));
    OR2B count_n1_0_i_o3 (.A(scalestate_0_dump_sustain_ctrl), .B(
        AND2_1_Y), .Y(N_11));
    
endmodule


module cal_load(
       cal_data,
       cal_para_out,
       top_code_0_cal_load,
       GLA
    );
input  [5:0] cal_data;
output [5:0] cal_para_out;
input  top_code_0_cal_load;
input  GLA;

    wire GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1E1 \cal_para_out[5]  (.D(cal_data[5]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[5]));
    GND GND_i_0 (.Y(GND_0));
    DFN1E1 \cal_para_out[1]  (.D(cal_data[1]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[1]));
    DFN1E1 \cal_para_out[4]  (.D(cal_data[4]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[4]));
    DFN1E1 \cal_para_out[3]  (.D(cal_data[3]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[3]));
    DFN1E1 \cal_para_out[0]  (.D(cal_data[0]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[0]));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    DFN1E1 \cal_para_out[2]  (.D(cal_data[2]), .CLK(GLA), .E(
        top_code_0_cal_load), .Q(cal_para_out[2]));
    
endmodule


module cal_div(
       cal_para_out,
       ddsclkout_c,
       cal_out_c,
       net_33,
       scanstate_0_calctrl
    );
input  [5:0] cal_para_out;
input  ddsclkout_c;
output cal_out_c;
input  net_33;
input  scanstate_0_calctrl;

    wire N_15, \count[1]_net_1 , \count[0]_net_1 , N_7, 
        \count[3]_net_1 , \DWACT_FINC_E[0] , clear_n4_NE_3, 
        clear_n4_4_i, clear_n4_5_i, clear_n4_NE_1, clear_n4_NE_2, 
        clear_n4_0_i, \count[2]_net_1 , clear_n4_3_i, cal_1_sqmuxa_1, 
        cal_RNO_net_1, N_37, \count_5[0] , \count_5[5] , I_24_0, 
        \count_5[4] , I_20_0, \count_5[3] , I_13_0, \count_5[2] , 
        I_9_0, \count_5[1] , I_5_0, \count[5]_net_1 , \count[4]_net_1 , 
        N_4, N_12, GND, VCC, GND_0, VCC_0;
    
    DFN1 \count[5]  (.D(\count_5[5] ), .CLK(ddsclkout_c), .Q(
        \count[5]_net_1 ));
    DFN1 \count[1]  (.D(\count_5[1] ), .CLK(ddsclkout_c), .Q(
        \count[1]_net_1 ));
    DFN1 \count[0]  (.D(\count_5[0] ), .CLK(ddsclkout_c), .Q(
        \count[0]_net_1 ));
    AND3 un3_count_I_16 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(\DWACT_FINC_E[0] ));
    NOR2B cal_RNO (.A(net_33), .B(N_37), .Y(cal_RNO_net_1));
    NOR3C \count_RNO[2]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(I_9_0), 
        .Y(\count_5[2] ));
    AOI1B \count_RNIQ24H1[1]  (.A(clear_n4_NE_3), .B(clear_n4_NE_2), 
        .C(scanstate_0_calctrl), .Y(cal_1_sqmuxa_1));
    NOR3C \count_RNICMJS[2]  (.A(clear_n4_4_i), .B(clear_n4_5_i), .C(
        clear_n4_NE_1), .Y(clear_n4_NE_3));
    XA1A \count_RNI2B9E[2]  (.A(\count[2]_net_1 ), .B(cal_para_out[2]), 
        .C(clear_n4_3_i), .Y(clear_n4_NE_1));
    VCC VCC_i (.Y(VCC));
    NOR3C \count_RNO[4]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(I_20_0), 
        .Y(\count_5[4] ));
    XNOR2 \count_RNIM957[5]  (.A(cal_para_out[5]), .B(\count[5]_net_1 )
        , .Y(clear_n4_5_i));
    XOR2 un3_count_I_5 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), .Y(
        I_5_0));
    NOR3C \count_RNO[3]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(I_13_0), 
        .Y(\count_5[3] ));
    NOR3C \count_RNO[5]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(I_24_0), 
        .Y(\count_5[5] ));
    NOR3C \count_RNO[1]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(I_5_0), 
        .Y(\count_5[1] ));
    XNOR2 \count_RNIK157[4]  (.A(cal_para_out[4]), .B(\count[4]_net_1 )
        , .Y(clear_n4_4_i));
    XOR2 un3_count_I_9 (.A(N_15), .B(\count[2]_net_1 ), .Y(I_9_0));
    DFN1 \count[2]  (.D(\count_5[2] ), .CLK(ddsclkout_c), .Q(
        \count[2]_net_1 ));
    XA1A \count_RNIQA8E[1]  (.A(\count[1]_net_1 ), .B(cal_para_out[1]), 
        .C(clear_n4_0_i), .Y(clear_n4_NE_2));
    XOR2 un3_count_I_24 (.A(N_4), .B(\count[5]_net_1 ), .Y(I_24_0));
    GND GND_i (.Y(GND));
    NOR2B un3_count_I_19 (.A(\count[3]_net_1 ), .B(\DWACT_FINC_E[0] ), 
        .Y(N_7));
    AND3 un3_count_I_12 (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(\count[2]_net_1 ), .Y(N_12));
    OR3C \count_RNO[0]  (.A(cal_1_sqmuxa_1), .B(net_33), .C(
        \count[0]_net_1 ), .Y(\count_5[0] ));
    NOR2B un3_count_I_8 (.A(\count[1]_net_1 ), .B(\count[0]_net_1 ), 
        .Y(N_15));
    DFN1 \count[3]  (.D(\count_5[3] ), .CLK(ddsclkout_c), .Q(
        \count[3]_net_1 ));
    AXOI7 cal_RNO_0 (.A(scanstate_0_calctrl), .B(cal_1_sqmuxa_1), .C(
        cal_out_c), .Y(N_37));
    XNOR2 \count_RNIC147[0]  (.A(cal_para_out[0]), .B(\count[0]_net_1 )
        , .Y(clear_n4_0_i));
    XOR2 un3_count_I_20 (.A(N_7), .B(\count[4]_net_1 ), .Y(I_20_0));
    DFN1 cal (.D(cal_RNO_net_1), .CLK(ddsclkout_c), .Q(cal_out_c));
    XNOR2 \count_RNIIP47[3]  (.A(cal_para_out[3]), .B(\count[3]_net_1 )
        , .Y(clear_n4_3_i));
    DFN1 \count[4]  (.D(\count_5[4] ), .CLK(ddsclkout_c), .Q(
        \count[4]_net_1 ));
    AND3 un3_count_I_23 (.A(\DWACT_FINC_E[0] ), .B(\count[3]_net_1 ), 
        .C(\count[4]_net_1 ), .Y(N_4));
    XOR2 un3_count_I_13 (.A(N_12), .B(\count[3]_net_1 ), .Y(I_13_0));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module CAL(
       cal_data,
       scanstate_0_calctrl,
       net_33,
       cal_out_c,
       ddsclkout_c,
       GLA,
       top_code_0_cal_load
    );
input  [5:0] cal_data;
input  scanstate_0_calctrl;
input  net_33;
output cal_out_c;
input  ddsclkout_c;
input  GLA;
input  top_code_0_cal_load;

    wire \cal_para_out[0] , \cal_para_out[1] , \cal_para_out[2] , 
        \cal_para_out[3] , \cal_para_out[4] , \cal_para_out[5] , GND, 
        VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    cal_load cal_load_0 (.cal_data({cal_data[5], cal_data[4], 
        cal_data[3], cal_data[2], cal_data[1], cal_data[0]}), 
        .cal_para_out({\cal_para_out[5] , \cal_para_out[4] , 
        \cal_para_out[3] , \cal_para_out[2] , \cal_para_out[1] , 
        \cal_para_out[0] }), .top_code_0_cal_load(top_code_0_cal_load), 
        .GLA(GLA));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    cal_div cal_div_0 (.cal_para_out({\cal_para_out[5] , 
        \cal_para_out[4] , \cal_para_out[3] , \cal_para_out[2] , 
        \cal_para_out[1] , \cal_para_out[0] }), .ddsclkout_c(
        ddsclkout_c), .cal_out_c(cal_out_c), .net_33(net_33), 
        .scanstate_0_calctrl(scanstate_0_calctrl));
    
endmodule


module qq_state_qq_state_0(
       i_1,
       i_2,
       GLA,
       Q1Q8_c,
       qq_state_0_stateover,
       Q3Q6_c,
       bri_dump_sw_0_reset_out_0
    );
input  [3:1] i_1;
input  [0:0] i_2;
input  GLA;
output Q1Q8_c;
output qq_state_0_stateover;
output Q3Q6_c;
input  bri_dump_sw_0_reset_out_0;

    wire \cs_RNO[2]_net_1 , cs4, N_89, N_88, \cs_RNO[3]_net_1 , N_86, 
        N_87, Q1Q8_Q2Q7_RNO_net_1, N_79, \cs[4]_net_1 , N_84, 
        \cs[3]_net_1 , \cs[1]_net_1 , \cs_RNO[1]_net_1 , 
        \cs_i[0]_net_1 , N_82, \cs_RNO[4]_net_1 , stateover_RNO_net_1, 
        GND, VCC, GND_0, VCC_0;
    
    AO1B stateover_RNO (.A(qq_state_0_stateover), .B(N_84), .C(cs4), 
        .Y(stateover_RNO_net_1));
    DFN1 \cs[2]  (.D(\cs_RNO[2]_net_1 ), .CLK(GLA), .Q(Q3Q6_c));
    NOR2B cs4_0_o3 (.A(bri_dump_sw_0_reset_out_0), .B(i_2[0]), .Y(cs4));
    GND GND_i_0 (.Y(GND_0));
    NOR2 \cs_RNO_1[3]  (.A(i_1[2]), .B(\cs[3]_net_1 ), .Y(N_87));
    NOR3A Q1Q8_Q2Q7_RNO (.A(cs4), .B(N_79), .C(\cs[4]_net_1 ), .Y(
        Q1Q8_Q2Q7_RNO_net_1));
    OA1C \cs_RNO_0[3]  (.A(\cs[3]_net_1 ), .B(i_1[3]), .C(Q3Q6_c), .Y(
        N_86));
    DFN1 \cs[3]  (.D(\cs_RNO[3]_net_1 ), .CLK(GLA), .Q(\cs[3]_net_1 ));
    NOR3A \cs_RNO[3]  (.A(cs4), .B(N_86), .C(N_87), .Y(
        \cs_RNO[3]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1 \cs[4]  (.D(\cs_RNO[4]_net_1 ), .CLK(GLA), .Q(\cs[4]_net_1 ));
    DFN1 stateover (.D(stateover_RNO_net_1), .CLK(GLA), .Q(
        qq_state_0_stateover));
    AOI1B \cs_RNO[1]  (.A(\cs_i[0]_net_1 ), .B(N_82), .C(cs4), .Y(
        \cs_RNO[1]_net_1 ));
    GND GND_i (.Y(GND));
    OR2A \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_1[1]), .Y(N_82));
    NOR2B \cs_RNI1E06[3]  (.A(i_1[3]), .B(\cs[3]_net_1 ), .Y(N_79));
    NOR2 \cs_RNO_1[2]  (.A(Q3Q6_c), .B(i_1[1]), .Y(N_88));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2A \cs_RNO[4]  (.A(cs4), .B(N_84), .Y(\cs_RNO[4]_net_1 ));
    DFN1 \cs[1]  (.D(\cs_RNO[1]_net_1 ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    DFN1 \cs_i[0]  (.D(cs4), .CLK(GLA), .Q(\cs_i[0]_net_1 ));
    DFN1 Q1Q8_Q2Q7 (.D(Q1Q8_Q2Q7_RNO_net_1), .CLK(GLA), .Q(Q1Q8_c));
    OA1C \cs_RNO_0[2]  (.A(Q3Q6_c), .B(i_1[2]), .C(\cs[1]_net_1 ), .Y(
        N_89));
    NOR3A \cs_RNO[2]  (.A(cs4), .B(N_89), .C(N_88), .Y(
        \cs_RNO[2]_net_1 ));
    NOR2 \cs_RNIGLBB[4]  (.A(\cs[4]_net_1 ), .B(N_79), .Y(N_84));
    
endmodule


module qq_coder_qq_coder_0(
       i_1,
       i_2,
       qq_para2,
       qq_para3,
       count_1,
       qq_para1,
       GLA,
       up,
       bri_dump_sw_0_reset_out_0
    );
output [3:1] i_1;
output [0:0] i_2;
input  [5:0] qq_para2;
input  [5:0] qq_para3;
input  [4:0] count_1;
input  [3:0] qq_para1;
input  GLA;
input  up;
input  bri_dump_sw_0_reset_out_0;

    wire \i_0_4[1] , \i_0_1[1] , \i_0_2[1] , \i_0_0[1] , 
        \un1_count_3_i_0[0] , \i_reg10_NE_3[0]_net_1 , 
        \i_reg10_2_i[0] , \i_reg10_1_i[0] , \i_reg10_NE_0[0]_net_1 , 
        \i_reg10_NE_2[0]_net_1 , \i_reg10_0_i[0] , 
        \un1_qq_para2_NE_2[0]_net_1 , \un1_qq_para2_0_i[0] , 
        \un1_qq_para2_NE_1[0]_net_1 , \un1_qq_para2_2_i[0] , 
        \un1_qq_para2_NE_0[0]_net_1 , \i_RNO[1]_net_1 , 
        \un1_qq_para2_i[0] , \i_reg10_NE_i_0[0] , \i_RNO[2]_net_1 , 
        \i_RNO[0]_net_1 , \i_RNO[3]_net_1 , GND, VCC, GND_0, VCC_0;
    
    XNOR2 \un1_qq_para2_2_0[0]  (.A(count_1[2]), .B(qq_para2[2]), .Y(
        \un1_qq_para2_2_i[0] ));
    XA1C \i_RNO_4[1]  (.A(qq_para1[1]), .B(count_1[1]), .C(count_1[4]), 
        .Y(\i_0_0[1] ));
    XA1A \i_reg10_NE_2[0]  (.A(qq_para3[3]), .B(count_1[3]), .C(
        \i_reg10_0_i[0] ), .Y(\i_reg10_NE_2[0]_net_1 ));
    DFN1 \i[3]  (.D(\i_RNO[3]_net_1 ), .CLK(GLA), .Q(i_1[3]));
    XNOR2 \i_reg10_1_0[0]  (.A(count_1[1]), .B(qq_para3[1]), .Y(
        \i_reg10_1_i[0] ));
    XA1C \i_reg10_NE_0[0]  (.A(qq_para3[4]), .B(count_1[4]), .C(
        qq_para3[5]), .Y(\i_reg10_NE_0[0]_net_1 ));
    XA1A \un1_qq_para2_NE_1[0]  (.A(qq_para2[1]), .B(count_1[1]), .C(
        \un1_qq_para2_2_i[0] ), .Y(\un1_qq_para2_NE_1[0]_net_1 ));
    DFN1 \i[0]  (.D(\i_RNO[0]_net_1 ), .CLK(GLA), .Q(i_2[0]));
    GND GND_i_0 (.Y(GND_0));
    DFN1 \i[2]  (.D(\i_RNO[2]_net_1 ), .CLK(GLA), .Q(i_1[2]));
    VCC VCC_i (.Y(VCC));
    XNOR2 \un1_qq_para2_0_0[0]  (.A(count_1[0]), .B(qq_para2[0]), .Y(
        \un1_qq_para2_0_i[0] ));
    NOR2B \i_RNO[0]  (.A(up), .B(bri_dump_sw_0_reset_out_0), .Y(
        \i_RNO[0]_net_1 ));
    NOR2B \i_RNO[3]  (.A(bri_dump_sw_0_reset_out_0), .B(
        \i_reg10_NE_i_0[0] ), .Y(\i_RNO[3]_net_1 ));
    NOR3B \i_RNO[1]  (.A(\i_0_4[1] ), .B(\un1_qq_para2_i[0] ), .C(
        \i_reg10_NE_i_0[0] ), .Y(\i_RNO[1]_net_1 ));
    XNOR2 \i_reg10_0_0[0]  (.A(count_1[0]), .B(qq_para3[0]), .Y(
        \i_reg10_0_i[0] ));
    GND GND_i (.Y(GND));
    XA1A \i_RNO_1[1]  (.A(qq_para1[2]), .B(count_1[2]), .C(
        \un1_count_3_i_0[0] ), .Y(\i_0_1[1] ));
    XA1C \un1_qq_para2_NE_0[0]  (.A(qq_para2[4]), .B(count_1[4]), .C(
        qq_para2[5]), .Y(\un1_qq_para2_NE_0[0]_net_1 ));
    NOR2B \i_reg10_NE[0]  (.A(\i_reg10_NE_3[0]_net_1 ), .B(
        \i_reg10_NE_2[0]_net_1 ), .Y(\i_reg10_NE_i_0[0] ));
    XNOR2 \i_reg10_2_0[0]  (.A(count_1[2]), .B(qq_para3[2]), .Y(
        \i_reg10_2_i[0] ));
    XA1A \i_RNO_2[1]  (.A(qq_para1[0]), .B(count_1[0]), .C(\i_0_0[1] ), 
        .Y(\i_0_2[1] ));
    DFN1 \i[1]  (.D(\i_RNO[1]_net_1 ), .CLK(GLA), .Q(i_1[1]));
    VCC VCC_i_0 (.Y(VCC_0));
    XNOR2 \i_RNO_3[1]  (.A(count_1[3]), .B(qq_para1[3]), .Y(
        \un1_count_3_i_0[0] ));
    NOR3C \i_reg10_NE_3[0]  (.A(\i_reg10_2_i[0] ), .B(\i_reg10_1_i[0] )
        , .C(\i_reg10_NE_0[0]_net_1 ), .Y(\i_reg10_NE_3[0]_net_1 ));
    NOR3C \i_RNO_0[1]  (.A(bri_dump_sw_0_reset_out_0), .B(\i_0_1[1] ), 
        .C(\i_0_2[1] ), .Y(\i_0_4[1] ));
    OR3C \un1_qq_para2_NE[0]  (.A(\un1_qq_para2_NE_1[0]_net_1 ), .B(
        \un1_qq_para2_NE_0[0]_net_1 ), .C(\un1_qq_para2_NE_2[0]_net_1 )
        , .Y(\un1_qq_para2_i[0] ));
    XA1A \un1_qq_para2_NE_2[0]  (.A(qq_para2[3]), .B(count_1[3]), .C(
        \un1_qq_para2_0_i[0] ), .Y(\un1_qq_para2_NE_2[0]_net_1 ));
    NOR3A \i_RNO[2]  (.A(bri_dump_sw_0_reset_out_0), .B(
        \un1_qq_para2_i[0] ), .C(\i_reg10_NE_i_0[0] ), .Y(
        \i_RNO[2]_net_1 ));
    
endmodule


module bri_timer(
       count,
       count_0,
       bri_dump_sw_0_reset_out,
       ddsclkout_c,
       bri_coder_0_half,
       pulse_start_c,
       clk_4f_en
    );
output [7:5] count;
output [4:0] count_0;
input  bri_dump_sw_0_reset_out;
input  ddsclkout_c;
input  bri_coder_0_half;
input  pulse_start_c;
input  clk_4f_en;

    wire clken_net_1, count_c2, count_c4, count_c5, count_n1, 
        \count_RNO[0]_net_1 , count_n2, count_n3, count_n4, count_n5, 
        count_n6, count_n7, GND, VCC, GND_0, VCC_0;
    
    XOR2 \count_RNO[6]  (.A(count[6]), .B(count_c5), .Y(count_n6));
    DFN1E1C0 \count[5]  (.D(count_n5), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count[5]));
    GND GND_i_0 (.Y(GND_0));
    XOR2 \count_RNO[1]  (.A(count_0[1]), .B(count_0[0]), .Y(count_n1));
    DFN1E1C0 \count[3]  (.D(count_n3), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count_0[3]));
    NOR3B clken (.A(clk_4f_en), .B(pulse_start_c), .C(bri_coder_0_half)
        , .Y(clken_net_1));
    DFN1C0 \count[0]  (.D(\count_RNO[0]_net_1 ), .CLK(ddsclkout_c), 
        .CLR(bri_dump_sw_0_reset_out), .Q(count_0[0]));
    XOR2 \count_RNO[3]  (.A(count_0[3]), .B(count_c2), .Y(count_n3));
    VCC VCC_i (.Y(VCC));
    XOR2 \count_RNO[5]  (.A(count[5]), .B(count_c4), .Y(count_n5));
    NOR3C \count_RNIUK31[0]  (.A(count_0[0]), .B(count_0[1]), .C(
        count_0[2]), .Y(count_c2));
    AX1C \count_RNO[7]  (.A(count_c5), .B(count[6]), .C(count[7]), .Y(
        count_n7));
    GND GND_i (.Y(GND));
    AX1C \count_RNO[2]  (.A(count_0[0]), .B(count_0[1]), .C(count_0[2])
        , .Y(count_n2));
    NOR3C \count_RNIN1S1[4]  (.A(count_c2), .B(count_0[3]), .C(
        count_0[4]), .Y(count_c4));
    VCC VCC_i_0 (.Y(VCC_0));
    AX1C \count_RNO[4]  (.A(count_c2), .B(count_0[3]), .C(count_0[4]), 
        .Y(count_n4));
    DFN1E1C0 \count[1]  (.D(count_n1), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count_0[1]));
    NOR2B \count_RNI5E82[5]  (.A(count[5]), .B(count_c4), .Y(count_c5));
    DFN1E1C0 \count[4]  (.D(count_n4), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count_0[4]));
    XOR2 \count_RNO[0]  (.A(count_0[0]), .B(clken_net_1), .Y(
        \count_RNO[0]_net_1 ));
    DFN1E1C0 \count[6]  (.D(count_n6), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count[6]));
    DFN1E1C0 \count[7]  (.D(count_n7), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count[7]));
    DFN1E1C0 \count[2]  (.D(count_n2), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clken_net_1), .Q(count_0[2]));
    
endmodule


module bri_coder(
       half_para,
       i_0,
       i_1,
       count_0,
       count,
       net_51,
       bri_dump_sw_0_phase_ctr,
       bri_dump_sw_0_reset_out,
       clk_4f_en,
       pulse_start_c,
       bri_dump_sw_0_reset_out_0,
       ddsclkout_c,
       bri_coder_0_half,
       PLUSE_0_bri_cycle
    );
input  [7:0] half_para;
output [3:1] i_0;
output [0:0] i_1;
input  [4:0] count_0;
input  [7:5] count;
input  net_51;
input  bri_dump_sw_0_phase_ctr;
input  bri_dump_sw_0_reset_out;
input  clk_4f_en;
input  pulse_start_c;
input  bri_dump_sw_0_reset_out_0;
input  ddsclkout_c;
output bri_coder_0_half;
output PLUSE_0_bri_cycle;

    wire un2lto7_3_net_1, un2lto7_0_net_1, un2lto7_2_net_1, 
        \DWACT_COMP0_E[1] , \DWACT_COMP0_E[2] , \DWACT_COMP0_E[0] , 
        N_17, N_16, N_15, N_12, N_14, N_13, N_11, N_8, N_9, N_10, 
        \ACT_LT3_E[3] , \ACT_LT3_E[4] , \ACT_LT3_E[5] , \ACT_LT3_E[0] , 
        \ACT_LT3_E[1] , \ACT_LT3_E[2] , \DWACT_BL_EQUAL_0_E[2] , 
        \DWACT_BL_EQUAL_0_E[1] , \DWACT_BL_EQUAL_0_E[0] , GND, VCC, 
        GND_0, VCC_0;
    
    OA1A half_0_I_31 (.A(N_12), .B(N_14), .C(N_13), .Y(N_17));
    OA1A half_0_I_27 (.A(half_para[3]), .B(count_0[3]), .C(N_9), .Y(
        N_13));
    DFN1E1C0 \i[2]  (.D(bri_dump_sw_0_phase_ctr), .CLK(ddsclkout_c), 
        .CLR(bri_dump_sw_0_reset_out), .E(clk_4f_en), .Q(i_0[2]));
    AOI1 bri_cycle (.A(un2lto7_3_net_1), .B(un2lto7_2_net_1), .C(
        bri_coder_0_half), .Y(PLUSE_0_bri_cycle));
    DFN1E1C0 \i[3]  (.D(net_51), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clk_4f_en), .Q(i_0[3]));
    OA1 half_0_I_32 (.A(N_17), .B(N_16), .C(N_15), .Y(
        \DWACT_COMP0_E[2] ));
    XNOR2 half_0_I_1 (.A(half_para[5]), .B(count[5]), .Y(
        \DWACT_BL_EQUAL_0_E[0] ));
    NOR2 un2lto7_2 (.A(count[6]), .B(count[7]), .Y(un2lto7_2_net_1));
    OR2A half_0_I_22 (.A(count_0[1]), .B(half_para[1]), .Y(N_8));
    VCC VCC_i (.Y(VCC));
    AO1C half_0_I_30 (.A(half_para[3]), .B(count_0[3]), .C(N_11), .Y(
        N_16));
    AND2A half_0_I_11 (.A(count[6]), .B(half_para[6]), .Y(
        \ACT_LT3_E[2] ));
    AND3 half_0_I_4 (.A(\DWACT_BL_EQUAL_0_E[2] ), .B(
        \DWACT_BL_EQUAL_0_E[1] ), .C(\DWACT_BL_EQUAL_0_E[0] ), .Y(
        \DWACT_COMP0_E[1] ));
    OR2A half_0_I_23 (.A(half_para[2]), .B(count_0[2]), .Y(N_9));
    AO1C half_0_I_28 (.A(half_para[2]), .B(count_0[2]), .C(N_8), .Y(
        N_14));
    AOI1A half_0_I_12 (.A(\ACT_LT3_E[0] ), .B(\ACT_LT3_E[1] ), .C(
        \ACT_LT3_E[2] ), .Y(\ACT_LT3_E[3] ));
    OR2A half_0_I_13 (.A(count[7]), .B(half_para[7]), .Y(
        \ACT_LT3_E[4] ));
    OR2A half_0_I_10 (.A(count[6]), .B(half_para[6]), .Y(
        \ACT_LT3_E[1] ));
    DFN1E1C0 \i[0]  (.D(pulse_start_c), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out_0), .E(clk_4f_en), .Q(i_1[0]));
    NOR2A half_0_I_24 (.A(count_0[0]), .B(half_para[0]), .Y(N_10));
    GND GND_i (.Y(GND));
    AO1C half_0_I_26 (.A(count_0[1]), .B(half_para[1]), .C(N_10), .Y(
        N_12));
    NOR2A half_0_I_9 (.A(count[5]), .B(half_para[5]), .Y(
        \ACT_LT3_E[0] ));
    AND2A half_0_I_14 (.A(count[7]), .B(half_para[7]), .Y(
        \ACT_LT3_E[5] ));
    OR2A half_0_I_25 (.A(count_0[4]), .B(half_para[4]), .Y(N_11));
    AOI1 un2lto7_0 (.A(count_0[2]), .B(count_0[1]), .C(count_0[3]), .Y(
        un2lto7_0_net_1));
    AO1 half_0_I_39 (.A(\DWACT_COMP0_E[1] ), .B(\DWACT_COMP0_E[2] ), 
        .C(\DWACT_COMP0_E[0] ), .Y(bri_coder_0_half));
    AOI1A half_0_I_15 (.A(\ACT_LT3_E[3] ), .B(\ACT_LT3_E[4] ), .C(
        \ACT_LT3_E[5] ), .Y(\DWACT_COMP0_E[0] ));
    NOR3A un2lto7_3 (.A(un2lto7_0_net_1), .B(count[5]), .C(count_0[4]), 
        .Y(un2lto7_3_net_1));
    XNOR2 half_0_I_3 (.A(half_para[7]), .B(count[7]), .Y(
        \DWACT_BL_EQUAL_0_E[2] ));
    OR2A half_0_I_29 (.A(half_para[4]), .B(count_0[4]), .Y(N_15));
    DFN1E1C0 \i[1]  (.D(bri_coder_0_half), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clk_4f_en), .Q(i_0[1]));
    VCC VCC_i_0 (.Y(VCC_0));
    XNOR2 half_0_I_2 (.A(half_para[6]), .B(count[6]), .Y(
        \DWACT_BL_EQUAL_0_E[1] ));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module qq_state_qq_state_0_1(
       i,
       i_0,
       GLA,
       Q2Q7_c,
       qq_state_1_stateover,
       Q4Q5_c,
       bri_dump_sw_0_reset_out_0
    );
input  [3:1] i;
input  [0:0] i_0;
input  GLA;
output Q2Q7_c;
output qq_state_1_stateover;
output Q4Q5_c;
input  bri_dump_sw_0_reset_out_0;

    wire N_77, cs4, N_89, N_88, N_71, N_86, N_87, N_65, N_79, 
        \cs[4]_net_1 , N_84, \cs[3]_net_1 , \cs[1]_net_1 , N_67, 
        \cs_i[0]_net_1 , N_82, N_73, N_34, GND, VCC, GND_0, VCC_0;
    
    AO1B stateover_RNO (.A(qq_state_1_stateover), .B(N_84), .C(cs4), 
        .Y(N_34));
    NOR2 \cs_RNIJLBB[4]  (.A(\cs[4]_net_1 ), .B(N_79), .Y(N_84));
    DFN1 \cs[2]  (.D(N_77), .CLK(GLA), .Q(Q4Q5_c));
    NOR2B cs4_0_o3 (.A(bri_dump_sw_0_reset_out_0), .B(i_0[0]), .Y(cs4));
    GND GND_i_0 (.Y(GND_0));
    NOR2 \cs_RNO_1[3]  (.A(i[2]), .B(\cs[3]_net_1 ), .Y(N_87));
    NOR3A Q1Q8_Q2Q7_RNO (.A(cs4), .B(N_79), .C(\cs[4]_net_1 ), .Y(N_65)
        );
    OA1C \cs_RNO_0[3]  (.A(\cs[3]_net_1 ), .B(i[3]), .C(Q4Q5_c), .Y(
        N_86));
    DFN1 \cs[3]  (.D(N_71), .CLK(GLA), .Q(\cs[3]_net_1 ));
    NOR3A \cs_RNO[3]  (.A(cs4), .B(N_86), .C(N_87), .Y(N_71));
    VCC VCC_i (.Y(VCC));
    DFN1 \cs[4]  (.D(N_73), .CLK(GLA), .Q(\cs[4]_net_1 ));
    DFN1 stateover (.D(N_34), .CLK(GLA), .Q(qq_state_1_stateover));
    AOI1B \cs_RNO[1]  (.A(\cs_i[0]_net_1 ), .B(N_82), .C(cs4), .Y(N_67)
        );
    GND GND_i (.Y(GND));
    NOR2B \cs_RNI3E06[3]  (.A(i[3]), .B(\cs[3]_net_1 ), .Y(N_79));
    OR2A \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i[1]), .Y(N_82));
    NOR2 \cs_RNO_1[2]  (.A(Q4Q5_c), .B(i[1]), .Y(N_88));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2A \cs_RNO[4]  (.A(cs4), .B(N_84), .Y(N_73));
    DFN1 \cs[1]  (.D(N_67), .CLK(GLA), .Q(\cs[1]_net_1 ));
    DFN1 \cs_i[0]  (.D(cs4), .CLK(GLA), .Q(\cs_i[0]_net_1 ));
    DFN1 Q1Q8_Q2Q7 (.D(N_65), .CLK(GLA), .Q(Q2Q7_c));
    OA1C \cs_RNO_0[2]  (.A(Q4Q5_c), .B(i[2]), .C(\cs[1]_net_1 ), .Y(
        N_89));
    NOR3A \cs_RNO[2]  (.A(cs4), .B(N_89), .C(N_88), .Y(N_77));
    
endmodule


module qq_timer_qq_timer_0(
       count_1,
       GLA,
       bri_dump_sw_0_reset_out_0,
       up,
       qq_state_0_stateover
    );
output [4:0] count_1;
input  GLA;
input  bri_dump_sw_0_reset_out_0;
input  up;
input  qq_state_0_stateover;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_15_i, GND, VCC, GND_0, VCC_0;
    
    NOR2B \count_RNI5TDG[2]  (.A(count_1[2]), .B(N_12), .Y(N_13));
    NOR2B \count_RNIDJUA[1]  (.A(count_1[1]), .B(count_1[0]), .Y(N_12));
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_1[0]), .B(count_1[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_1[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_1[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count_1[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    AX1E \count_RNO_0[4]  (.A(N_13), .B(count_1[3]), .C(count_1[4]), 
        .Y(N_15_i));
    XA1B \count_RNO[2]  (.A(N_12), .B(count_1[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(qq_state_0_stateover), .B(up), .C(
        bri_dump_sw_0_reset_out_0), .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \count_RNO[4]  (.A(count_0_sqmuxa_net_1), .B(N_15_i), .Y(N_11)
        );
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_1[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_1[4]));
    NOR2 \count_RNO[0]  (.A(count_1[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_1[2]));
    
endmodule


module qq_timer_qq_timer_0_1(
       count,
       GLA,
       bri_dump_sw_0_reset_out_0,
       down,
       qq_state_1_stateover
    );
output [4:0] count;
input  GLA;
input  bri_dump_sw_0_reset_out_0;
input  down;
input  qq_state_1_stateover;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_15_i, GND, VCC, GND_0, VCC_0;
    
    NOR2B \count_RNIFJUA[1]  (.A(count[1]), .B(count[0]), .Y(N_12));
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count[0]), .B(count[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    AX1E \count_RNO_0[4]  (.A(N_13), .B(count[3]), .C(count[4]), .Y(
        N_15_i));
    XA1B \count_RNO[2]  (.A(N_12), .B(count[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    NOR2B \count_RNI8TDG[2]  (.A(count[2]), .B(N_12), .Y(N_13));
    OR3C count_0_sqmuxa (.A(qq_state_1_stateover), .B(down), .C(
        bri_dump_sw_0_reset_out_0), .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \count_RNO[4]  (.A(count_0_sqmuxa_net_1), .B(N_15_i), .Y(N_11)
        );
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count[4]));
    NOR2 \count_RNO[0]  (.A(count[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count[2]));
    
endmodule


module qq_coder_qq_coder_0_1(
       i,
       i_0,
       qq_para2,
       qq_para3,
       count,
       qq_para1,
       GLA,
       down,
       bri_dump_sw_0_reset_out_0
    );
output [3:1] i;
output [0:0] i_0;
input  [5:0] qq_para2;
input  [5:0] qq_para3;
input  [4:0] count;
input  [3:0] qq_para1;
input  GLA;
input  down;
input  bri_dump_sw_0_reset_out_0;

    wire \i_0_4[1] , \i_0_1[1] , \i_0_2[1] , \i_0_0[1] , 
        \un1_count_3_i_0[0] , \i_reg10_NE_3[0]_net_1 , 
        \i_reg10_2_i[0] , \i_reg10_1_i[0] , \i_reg10_NE_0[0]_net_1 , 
        \i_reg10_NE_2[0]_net_1 , \i_reg10_0_i[0] , 
        \un1_qq_para2_NE_2[0]_net_1 , \un1_qq_para2_0_i[0] , 
        \un1_qq_para2_NE_1[0]_net_1 , \un1_qq_para2_2_i[0] , 
        \un1_qq_para2_NE_0[0]_net_1 , N_8, \un1_qq_para2_i[0] , 
        \i_reg10_NE_i_0[0] , N_9, N_7, N_10, GND, VCC, GND_0, VCC_0;
    
    XNOR2 \un1_qq_para2_2_0[0]  (.A(count[2]), .B(qq_para2[2]), .Y(
        \un1_qq_para2_2_i[0] ));
    XA1C \i_RNO_4[1]  (.A(qq_para1[1]), .B(count[1]), .C(count[4]), .Y(
        \i_0_0[1] ));
    XA1A \i_reg10_NE_2[0]  (.A(qq_para3[3]), .B(count[3]), .C(
        \i_reg10_0_i[0] ), .Y(\i_reg10_NE_2[0]_net_1 ));
    DFN1 \i[3]  (.D(N_10), .CLK(GLA), .Q(i[3]));
    XNOR2 \i_reg10_1_0[0]  (.A(count[1]), .B(qq_para3[1]), .Y(
        \i_reg10_1_i[0] ));
    XA1C \i_reg10_NE_0[0]  (.A(qq_para3[4]), .B(count[4]), .C(
        qq_para3[5]), .Y(\i_reg10_NE_0[0]_net_1 ));
    XA1A \un1_qq_para2_NE_1[0]  (.A(qq_para2[1]), .B(count[1]), .C(
        \un1_qq_para2_2_i[0] ), .Y(\un1_qq_para2_NE_1[0]_net_1 ));
    DFN1 \i[0]  (.D(N_7), .CLK(GLA), .Q(i_0[0]));
    GND GND_i_0 (.Y(GND_0));
    DFN1 \i[2]  (.D(N_9), .CLK(GLA), .Q(i[2]));
    VCC VCC_i (.Y(VCC));
    XNOR2 \un1_qq_para2_0_0[0]  (.A(count[0]), .B(qq_para2[0]), .Y(
        \un1_qq_para2_0_i[0] ));
    NOR2B \i_RNO[0]  (.A(down), .B(bri_dump_sw_0_reset_out_0), .Y(N_7));
    NOR2B \i_RNO[3]  (.A(bri_dump_sw_0_reset_out_0), .B(
        \i_reg10_NE_i_0[0] ), .Y(N_10));
    NOR3B \i_RNO[1]  (.A(\i_0_4[1] ), .B(\un1_qq_para2_i[0] ), .C(
        \i_reg10_NE_i_0[0] ), .Y(N_8));
    XNOR2 \i_reg10_0_0[0]  (.A(count[0]), .B(qq_para3[0]), .Y(
        \i_reg10_0_i[0] ));
    GND GND_i (.Y(GND));
    XA1A \i_RNO_1[1]  (.A(qq_para1[2]), .B(count[2]), .C(
        \un1_count_3_i_0[0] ), .Y(\i_0_1[1] ));
    XA1C \un1_qq_para2_NE_0[0]  (.A(qq_para2[4]), .B(count[4]), .C(
        qq_para2[5]), .Y(\un1_qq_para2_NE_0[0]_net_1 ));
    NOR2B \i_reg10_NE[0]  (.A(\i_reg10_NE_3[0]_net_1 ), .B(
        \i_reg10_NE_2[0]_net_1 ), .Y(\i_reg10_NE_i_0[0] ));
    XNOR2 \i_reg10_2_0[0]  (.A(count[2]), .B(qq_para3[2]), .Y(
        \i_reg10_2_i[0] ));
    XA1A \i_RNO_2[1]  (.A(qq_para1[0]), .B(count[0]), .C(\i_0_0[1] ), 
        .Y(\i_0_2[1] ));
    DFN1 \i[1]  (.D(N_8), .CLK(GLA), .Q(i[1]));
    VCC VCC_i_0 (.Y(VCC_0));
    XNOR2 \i_RNO_3[1]  (.A(count[3]), .B(qq_para1[3]), .Y(
        \un1_count_3_i_0[0] ));
    NOR3C \i_reg10_NE_3[0]  (.A(\i_reg10_2_i[0] ), .B(\i_reg10_1_i[0] )
        , .C(\i_reg10_NE_0[0]_net_1 ), .Y(\i_reg10_NE_3[0]_net_1 ));
    NOR3C \i_RNO_0[1]  (.A(bri_dump_sw_0_reset_out_0), .B(\i_0_1[1] ), 
        .C(\i_0_2[1] ), .Y(\i_0_4[1] ));
    OR3C \un1_qq_para2_NE[0]  (.A(\un1_qq_para2_NE_1[0]_net_1 ), .B(
        \un1_qq_para2_NE_0[0]_net_1 ), .C(\un1_qq_para2_NE_2[0]_net_1 )
        , .Y(\un1_qq_para2_i[0] ));
    XA1A \un1_qq_para2_NE_2[0]  (.A(qq_para2[3]), .B(count[3]), .C(
        \un1_qq_para2_0_i[0] ), .Y(\un1_qq_para2_NE_2[0]_net_1 ));
    NOR3A \i_RNO[2]  (.A(bri_dump_sw_0_reset_out_0), .B(
        \un1_qq_para2_i[0] ), .C(\i_reg10_NE_i_0[0] ), .Y(N_9));
    
endmodule


module bri_state(
       i_1,
       i_0,
       down,
       ddsclkout_c,
       up,
       bri_dump_sw_0_reset_out_0,
       clk_4f_en
    );
input  [0:0] i_1;
input  [3:1] i_0;
output down;
input  ddsclkout_c;
output up;
input  bri_dump_sw_0_reset_out_0;
input  clk_4f_en;

    wire csse_1_0_1, N_140, csse_1_0_0, \cs[2]_net_1 , csse_1_0_a4_1_0, 
        csse_1_0_a4_2_9, csse_1_0_a4_2_6, csse_1_0_a4_2_5, 
        csse_1_0_a4_2_7, csse_1_0_a4_2_4, \cs[3]_net_1 , 
        csse_1_0_a4_2_2, \cs[7]_net_1 , \cs[6]_net_1 , \cs[5]_net_1 , 
        \cs[4]_net_1 , \cs[8]_net_1 , \cs[11]_net_1 , \cs[12]_net_1 , 
        down32_0_o4_0, N_174, csse_9_0_a4_0_0, \cs[9]_net_1 , N_138, 
        csse_3_0_a4_0_0, \cs[1]_net_1 , csse_0_0_a4_0_0, \cs[0]_net_1 , 
        N_141, N_173, \cs_ns_e[2] , N_176, down30, N_171, en_net_1, 
        \cs_ns_e[0] , N_172, \cs[10]_net_1 , \cs_RNO[13]_net_1 , 
        \cs[13]_net_1 , \cs_RNO[12]_net_1 , \cs_RNO[11]_net_1 , 
        \cs_ns_e[10] , \cs_RNO[9]_net_1 , \cs_ns_e[8] , 
        \cs_RNO[7]_net_1 , \cs_RNO[6]_net_1 , \cs_RNO[5]_net_1 , 
        \cs_ns_e[4] , \cs_RNO_0[3] , \cs_ns_e[1] , down32, GND, VCC, 
        GND_0, VCC_0;
    
    DFN1E1C0 up_inst_1 (.D(down30), .CLK(ddsclkout_c), .CLR(en_net_1), 
        .E(clk_4f_en), .Q(up));
    OA1 \cs_RNI83HA[1]  (.A(N_172), .B(\cs[1]_net_1 ), .C(i_0[2]), .Y(
        N_173));
    OR3 up_RNO (.A(N_171), .B(\cs[2]_net_1 ), .C(N_140), .Y(down30));
    MX2 \cs_RNO[13]  (.A(\cs[13]_net_1 ), .B(\cs[12]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[13]_net_1 ));
    OR2 \cs_RNINU1L[1]  (.A(down32_0_o4_0), .B(N_173), .Y(N_141));
    MX2 \cs_RNO[10]  (.A(\cs[10]_net_1 ), .B(csse_9_0_a4_0_0), .S(
        clk_4f_en), .Y(\cs_ns_e[10] ));
    DFN1C0 \cs[6]  (.D(\cs_RNO[6]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[6]_net_1 ));
    NOR2 \cs_RNO_8[2]  (.A(\cs[8]_net_1 ), .B(i_0[3]), .Y(
        csse_1_0_a4_2_4));
    MX2 \cs_RNO[11]  (.A(\cs[11]_net_1 ), .B(\cs[10]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[11]_net_1 ));
    AO1A \cs_RNI298C[13]  (.A(N_138), .B(\cs[9]_net_1 ), .C(
        \cs[13]_net_1 ), .Y(N_140));
    DFN1E1C0 down_inst_1 (.D(down32), .CLK(ddsclkout_c), .CLR(en_net_1)
        , .E(clk_4f_en), .Q(down));
    NOR3A \cs_RNO_3[2]  (.A(csse_1_0_a4_2_2), .B(\cs[7]_net_1 ), .C(
        \cs[6]_net_1 ), .Y(csse_1_0_a4_2_6));
    NOR2A \cs_RNIKJ85[0]  (.A(\cs[0]_net_1 ), .B(i_0[3]), .Y(N_172));
    DFN1C0 \cs[12]  (.D(\cs_RNO[12]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[12]_net_1 ));
    AOI1B \cs_RNO_2[2]  (.A(clk_4f_en), .B(N_140), .C(csse_1_0_0), .Y(
        csse_1_0_1));
    NOR2A \cs_RNO[0]  (.A(\cs[0]_net_1 ), .B(clk_4f_en), .Y(
        \cs_ns_e[0] ));
    VCC VCC_i (.Y(VCC));
    DFN1C0 \cs[3]  (.D(\cs_RNO_0[3] ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[3]_net_1 ));
    MX2 \cs_RNO[7]  (.A(\cs[7]_net_1 ), .B(\cs[6]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[7]_net_1 ));
    MX2 \cs_RNO[1]  (.A(\cs[1]_net_1 ), .B(csse_0_0_a4_0_0), .S(
        clk_4f_en), .Y(\cs_ns_e[1] ));
    MX2 \cs_RNO[9]  (.A(\cs[9]_net_1 ), .B(\cs[8]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[9]_net_1 ));
    DFN1C0 \cs[5]  (.D(\cs_RNO[5]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[5]_net_1 ));
    MX2 \cs_RNO[8]  (.A(\cs[8]_net_1 ), .B(N_141), .S(clk_4f_en), .Y(
        \cs_ns_e[8] ));
    DFN1C0 \cs[11]  (.D(\cs_RNO[11]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[11]_net_1 ));
    DFN1C0 \cs[13]  (.D(\cs_RNO[13]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[13]_net_1 ));
    DFN1C0 \cs[2]  (.D(\cs_ns_e[2] ), .CLK(ddsclkout_c), .CLR(en_net_1)
        , .Q(\cs[2]_net_1 ));
    NOR2B en (.A(bri_dump_sw_0_reset_out_0), .B(i_1[0]), .Y(en_net_1));
    MX2 \cs_RNO[12]  (.A(\cs[12]_net_1 ), .B(\cs[11]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[12]_net_1 ));
    DFN1P0 \cs[0]  (.D(\cs_ns_e[0] ), .CLK(ddsclkout_c), .PRE(en_net_1)
        , .Q(\cs[0]_net_1 ));
    NOR2 \cs_RNO_7[2]  (.A(\cs[11]_net_1 ), .B(\cs[12]_net_1 ), .Y(
        csse_1_0_a4_2_2));
    GND GND_i (.Y(GND));
    OR2 down_RNO (.A(\cs[8]_net_1 ), .B(N_141), .Y(down32));
    NOR2B \cs_RNO_0[10]  (.A(\cs[9]_net_1 ), .B(N_138), .Y(
        csse_9_0_a4_0_0));
    NOR2A \cs_RNO_9[2]  (.A(\cs[1]_net_1 ), .B(i_0[2]), .Y(
        csse_1_0_a4_1_0));
    NOR3A \cs_RNO_5[2]  (.A(csse_1_0_a4_2_4), .B(\cs[3]_net_1 ), .C(
        \cs[2]_net_1 ), .Y(csse_1_0_a4_2_7));
    OA1 \cs_RNIEJB7[3]  (.A(i_0[1]), .B(i_0[2]), .C(\cs[3]_net_1 ), .Y(
        N_174));
    DFN1C0 \cs[10]  (.D(\cs_ns_e[10] ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[10]_net_1 ));
    AO1C \cs_RNO[2]  (.A(N_176), .B(csse_1_0_a4_2_9), .C(csse_1_0_1), 
        .Y(\cs_ns_e[2] ));
    OR2A \cs_RNO_0[2]  (.A(clk_4f_en), .B(\cs[10]_net_1 ), .Y(N_176));
    MX2C \cs_RNO_6[2]  (.A(\cs[2]_net_1 ), .B(csse_1_0_a4_1_0), .S(
        clk_4f_en), .Y(csse_1_0_0));
    MX2 \cs_RNO[4]  (.A(\cs[4]_net_1 ), .B(csse_3_0_a4_0_0), .S(
        clk_4f_en), .Y(\cs_ns_e[4] ));
    DFN1C0 \cs[9]  (.D(\cs_RNO[9]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[9]_net_1 ));
    DFN1C0 \cs[8]  (.D(\cs_ns_e[8] ), .CLK(ddsclkout_c), .CLR(en_net_1)
        , .Q(\cs[8]_net_1 ));
    MX2 \cs_RNO[6]  (.A(\cs[6]_net_1 ), .B(\cs[5]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[6]_net_1 ));
    NOR2A csse_9_0_o2 (.A(i_0[2]), .B(i_0[1]), .Y(N_138));
    NOR3C \cs_RNO_1[2]  (.A(csse_1_0_a4_2_6), .B(csse_1_0_a4_2_5), .C(
        csse_1_0_a4_2_7), .Y(csse_1_0_a4_2_9));
    OA1B up_RNO_0 (.A(N_172), .B(\cs[1]_net_1 ), .C(i_0[2]), .Y(N_171));
    NOR3 \cs_RNO_4[2]  (.A(\cs[5]_net_1 ), .B(\cs[4]_net_1 ), .C(
        i_0[2]), .Y(csse_1_0_a4_2_5));
    OR2 \cs_RNIFRGA[7]  (.A(\cs[7]_net_1 ), .B(N_174), .Y(
        down32_0_o4_0));
    MX2 \cs_RNO[3]  (.A(\cs[3]_net_1 ), .B(\cs[2]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO_0[3] ));
    DFN1C0 \cs[1]  (.D(\cs_ns_e[1] ), .CLK(ddsclkout_c), .CLR(en_net_1)
        , .Q(\cs[1]_net_1 ));
    MX2 \cs_RNO[5]  (.A(\cs[5]_net_1 ), .B(\cs[4]_net_1 ), .S(
        clk_4f_en), .Y(\cs_RNO[5]_net_1 ));
    DFN1C0 \cs[4]  (.D(\cs_ns_e[4] ), .CLK(ddsclkout_c), .CLR(en_net_1)
        , .Q(\cs[4]_net_1 ));
    DFN1C0 \cs[7]  (.D(\cs_RNO[7]_net_1 ), .CLK(ddsclkout_c), .CLR(
        en_net_1), .Q(\cs[7]_net_1 ));
    NOR2B \cs_RNO_0[1]  (.A(\cs[0]_net_1 ), .B(i_0[3]), .Y(
        csse_0_0_a4_0_0));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR3A \cs_RNO_0[4]  (.A(\cs[3]_net_1 ), .B(i_0[1]), .C(i_0[2]), .Y(
        csse_3_0_a4_0_0));
    
endmodule


module bri_qq_load(
       halfdata,
       half_para,
       qq_para1,
       qq_para2,
       bri_datain,
       qq_para3,
       top_code_0_bridge_load_0,
       top_code_0_bridge_load,
       GLA
    );
input  [7:0] halfdata;
output [7:0] half_para;
output [3:0] qq_para1;
output [5:0] qq_para2;
input  [15:0] bri_datain;
output [5:0] qq_para3;
input  top_code_0_bridge_load_0;
input  top_code_0_bridge_load;
input  GLA;

    wire GND, VCC, GND_0, VCC_0;
    
    DFN1E1 \qq_para1[0]  (.D(bri_datain[0]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para1[0]));
    DFN1E1 \half_para[2]  (.D(halfdata[2]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[2]));
    DFN1E1 \qq_para2[1]  (.D(bri_datain[5]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para2[1]));
    DFN1E1 \half_para[4]  (.D(halfdata[4]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[4]));
    DFN1E1 \qq_para3[2]  (.D(bri_datain[12]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[2]));
    DFN1E1 \half_para[6]  (.D(halfdata[6]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[6]));
    DFN1E1 \qq_para3[4]  (.D(bri_datain[14]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[4]));
    DFN1E1 \half_para[1]  (.D(halfdata[1]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[1]));
    GND GND_i_0 (.Y(GND_0));
    DFN1E1 \qq_para1[3]  (.D(bri_datain[3]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para1[3]));
    VCC VCC_i (.Y(VCC));
    DFN1E1 \qq_para3[0]  (.D(bri_datain[10]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[0]));
    DFN1E1 \qq_para1[1]  (.D(bri_datain[1]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para1[1]));
    DFN1E1 \qq_para3[1]  (.D(bri_datain[11]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[1]));
    DFN1E1 \qq_para2[3]  (.D(bri_datain[7]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para2[3]));
    DFN1E1 \qq_para2[0]  (.D(bri_datain[4]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para2[0]));
    GND GND_i (.Y(GND));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1E1 \half_para[5]  (.D(halfdata[5]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[5]));
    DFN1E1 \qq_para2[4]  (.D(bri_datain[8]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para2[4]));
    DFN1E1 \half_para[3]  (.D(halfdata[3]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[3]));
    DFN1E1 \qq_para3[3]  (.D(bri_datain[13]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[3]));
    DFN1E1 \qq_para2[2]  (.D(bri_datain[6]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para2[2]));
    DFN1E1 \qq_para3[5]  (.D(bri_datain[15]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para3[5]));
    DFN1E1 \qq_para2[5]  (.D(bri_datain[9]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(qq_para2[5]));
    DFN1E1 \qq_para1[2]  (.D(bri_datain[2]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(qq_para1[2]));
    DFN1E1 \half_para[0]  (.D(halfdata[0]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[0]));
    DFN1E1 \half_para[7]  (.D(halfdata[7]), .CLK(GLA), .E(
        top_code_0_bridge_load_0), .Q(half_para[7]));
    
endmodule


module PLUSE(
       bri_datain,
       halfdata,
       top_code_0_bridge_load,
       top_code_0_bridge_load_0,
       Q4Q5_c,
       Q2Q7_c,
       PLUSE_0_bri_cycle,
       bri_dump_sw_0_phase_ctr,
       net_51,
       clk_4f_en,
       pulse_start_c,
       ddsclkout_c,
       bri_dump_sw_0_reset_out,
       bri_dump_sw_0_reset_out_0,
       Q3Q6_c,
       Q1Q8_c,
       GLA
    );
input  [15:0] bri_datain;
input  [7:0] halfdata;
input  top_code_0_bridge_load;
input  top_code_0_bridge_load_0;
output Q4Q5_c;
output Q2Q7_c;
output PLUSE_0_bri_cycle;
input  bri_dump_sw_0_phase_ctr;
input  net_51;
input  clk_4f_en;
input  pulse_start_c;
input  ddsclkout_c;
input  bri_dump_sw_0_reset_out;
input  bri_dump_sw_0_reset_out_0;
output Q3Q6_c;
output Q1Q8_c;
input  GLA;

    wire \i_1[1] , \i_1[2] , \i_1[3] , \i_2[0] , qq_state_0_stateover, 
        \qq_para2[0] , \qq_para2[1] , \qq_para2[2] , \qq_para2[3] , 
        \qq_para2[4] , \qq_para2[5] , \qq_para3[0] , \qq_para3[1] , 
        \qq_para3[2] , \qq_para3[3] , \qq_para3[4] , \qq_para3[5] , 
        \count_1[0] , \count_1[1] , \count_1[2] , \count_1[3] , 
        \count_1[4] , \qq_para1[0] , \qq_para1[1] , \qq_para1[2] , 
        \qq_para1[3] , up, \count[5] , \count[6] , \count[7] , 
        \count_0[0] , \count_0[1] , \count_0[2] , \count_0[3] , 
        \count_0[4] , bri_coder_0_half, \half_para[0] , \half_para[1] , 
        \half_para[2] , \half_para[3] , \half_para[4] , \half_para[5] , 
        \half_para[6] , \half_para[7] , \i_0[1] , \i_0[2] , \i_0[3] , 
        \i_1[0] , \i[1] , \i[2] , \i[3] , \i_0[0] , 
        qq_state_1_stateover, \count[0] , \count[1] , \count[2] , 
        \count[3] , \count[4] , down, GND, VCC, GND_0, VCC_0;
    
    qq_state_qq_state_0 qq_state_0 (.i_1({\i_1[3] , \i_1[2] , \i_1[1] })
        , .i_2({\i_2[0] }), .GLA(GLA), .Q1Q8_c(Q1Q8_c), 
        .qq_state_0_stateover(qq_state_0_stateover), .Q3Q6_c(Q3Q6_c), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0));
    qq_coder_qq_coder_0 qq_coder_0 (.i_1({\i_1[3] , \i_1[2] , \i_1[1] })
        , .i_2({\i_2[0] }), .qq_para2({\qq_para2[5] , \qq_para2[4] , 
        \qq_para2[3] , \qq_para2[2] , \qq_para2[1] , \qq_para2[0] }), 
        .qq_para3({\qq_para3[5] , \qq_para3[4] , \qq_para3[3] , 
        \qq_para3[2] , \qq_para3[1] , \qq_para3[0] }), .count_1({
        \count_1[4] , \count_1[3] , \count_1[2] , \count_1[1] , 
        \count_1[0] }), .qq_para1({\qq_para1[3] , \qq_para1[2] , 
        \qq_para1[1] , \qq_para1[0] }), .GLA(GLA), .up(up), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0));
    bri_timer bri_timer_0 (.count({\count[7] , \count[6] , \count[5] })
        , .count_0({\count_0[4] , \count_0[3] , \count_0[2] , 
        \count_0[1] , \count_0[0] }), .bri_dump_sw_0_reset_out(
        bri_dump_sw_0_reset_out), .ddsclkout_c(ddsclkout_c), 
        .bri_coder_0_half(bri_coder_0_half), .pulse_start_c(
        pulse_start_c), .clk_4f_en(clk_4f_en));
    bri_coder bri_coder_0 (.half_para({\half_para[7] , \half_para[6] , 
        \half_para[5] , \half_para[4] , \half_para[3] , \half_para[2] , 
        \half_para[1] , \half_para[0] }), .i_0({\i_0[3] , \i_0[2] , 
        \i_0[1] }), .i_1({\i_1[0] }), .count_0({\count_0[4] , 
        \count_0[3] , \count_0[2] , \count_0[1] , \count_0[0] }), 
        .count({\count[7] , \count[6] , \count[5] }), .net_51(net_51), 
        .bri_dump_sw_0_phase_ctr(bri_dump_sw_0_phase_ctr), 
        .bri_dump_sw_0_reset_out(bri_dump_sw_0_reset_out), .clk_4f_en(
        clk_4f_en), .pulse_start_c(pulse_start_c), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), 
        .ddsclkout_c(ddsclkout_c), .bri_coder_0_half(bri_coder_0_half), 
        .PLUSE_0_bri_cycle(PLUSE_0_bri_cycle));
    qq_state_qq_state_0_1 qq_state_1 (.i({\i[3] , \i[2] , \i[1] }), 
        .i_0({\i_0[0] }), .GLA(GLA), .Q2Q7_c(Q2Q7_c), 
        .qq_state_1_stateover(qq_state_1_stateover), .Q4Q5_c(Q4Q5_c), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0));
    VCC VCC_i_0 (.Y(VCC_0));
    qq_timer_qq_timer_0 qq_timer_0 (.count_1({\count_1[4] , 
        \count_1[3] , \count_1[2] , \count_1[1] , \count_1[0] }), .GLA(
        GLA), .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), 
        .up(up), .qq_state_0_stateover(qq_state_0_stateover));
    VCC VCC_i (.Y(VCC));
    qq_timer_qq_timer_0_1 qq_timer_1 (.count({\count[4] , \count[3] , 
        \count[2] , \count[1] , \count[0] }), .GLA(GLA), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), .down(
        down), .qq_state_1_stateover(qq_state_1_stateover));
    qq_coder_qq_coder_0_1 qq_coder_1 (.i({\i[3] , \i[2] , \i[1] }), 
        .i_0({\i_0[0] }), .qq_para2({\qq_para2[5] , \qq_para2[4] , 
        \qq_para2[3] , \qq_para2[2] , \qq_para2[1] , \qq_para2[0] }), 
        .qq_para3({\qq_para3[5] , \qq_para3[4] , \qq_para3[3] , 
        \qq_para3[2] , \qq_para3[1] , \qq_para3[0] }), .count({
        \count[4] , \count[3] , \count[2] , \count[1] , \count[0] }), 
        .qq_para1({\qq_para1[3] , \qq_para1[2] , \qq_para1[1] , 
        \qq_para1[0] }), .GLA(GLA), .down(down), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    bri_state bri_state_0 (.i_1({\i_1[0] }), .i_0({\i_0[3] , \i_0[2] , 
        \i_0[1] }), .down(down), .ddsclkout_c(ddsclkout_c), .up(up), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), 
        .clk_4f_en(clk_4f_en));
    bri_qq_load bri_qq_load_0 (.halfdata({halfdata[7], halfdata[6], 
        halfdata[5], halfdata[4], halfdata[3], halfdata[2], 
        halfdata[1], halfdata[0]}), .half_para({\half_para[7] , 
        \half_para[6] , \half_para[5] , \half_para[4] , \half_para[3] , 
        \half_para[2] , \half_para[1] , \half_para[0] }), .qq_para1({
        \qq_para1[3] , \qq_para1[2] , \qq_para1[1] , \qq_para1[0] }), 
        .qq_para2({\qq_para2[5] , \qq_para2[4] , \qq_para2[3] , 
        \qq_para2[2] , \qq_para2[1] , \qq_para2[0] }), .bri_datain({
        bri_datain[15], bri_datain[14], bri_datain[13], bri_datain[12], 
        bri_datain[11], bri_datain[10], bri_datain[9], bri_datain[8], 
        bri_datain[7], bri_datain[6], bri_datain[5], bri_datain[4], 
        bri_datain[3], bri_datain[2], bri_datain[1], bri_datain[0]}), 
        .qq_para3({\qq_para3[5] , \qq_para3[4] , \qq_para3[3] , 
        \qq_para3[2] , \qq_para3[1] , \qq_para3[0] }), 
        .top_code_0_bridge_load_0(top_code_0_bridge_load_0), 
        .top_code_0_bridge_load(top_code_0_bridge_load), .GLA(GLA));
    
endmodule


module state_1ms(
       state_1ms_data,
       timecount_0,
       state_1ms_lc,
       GLA,
       state_1ms_0_reset_out,
       top_code_0_state_1ms_rst_n,
       top_code_0_state_1ms_load,
       state_1ms_0_bri_cycle,
       state_1ms_0_pluse_start,
       state_1ms_0_rt_sw,
       state_1ms_0_soft_dump,
       state_1ms_0_dump_start,
       top_code_0_state_1ms_rst_n_0,
       timer_top_0_clk_en_st1ms
    );
input  [15:0] state_1ms_data;
output [19:0] timecount_0;
input  [3:0] state_1ms_lc;
input  GLA;
output state_1ms_0_reset_out;
input  top_code_0_state_1ms_rst_n;
input  top_code_0_state_1ms_load;
output state_1ms_0_bri_cycle;
output state_1ms_0_pluse_start;
output state_1ms_0_rt_sw;
output state_1ms_0_soft_dump;
output state_1ms_0_dump_start;
input  top_code_0_state_1ms_rst_n_0;
input  timer_top_0_clk_en_st1ms;

    wire \timecount_8_iv_2[2] , \CS[7]_net_1 , \S_DUMPTIME[2]_net_1 , 
        \timecount_RNO_6[2]_net_1 , \timecount_8_iv_1[2] , 
        \CS[4]_net_1 , \PLUSECYCLE[2]_net_1 , 
        \timecount_RNO_5[2]_net_1 , \timecount_8_iv_0[2] , 
        \CS[6]_net_1 , \M_DUMPTIME[2]_net_1 , \CS_i[0]_net_1 , 
        \timecount_8_iv_2[5] , \S_DUMPTIME[5]_net_1 , 
        \timecount_RNO_6[5]_net_1 , \timecount_8_iv_1[5] , 
        \PLUSECYCLE[5]_net_1 , \timecount_RNO_5[5]_net_1 , 
        \timecount_8_iv_0[5] , \M_DUMPTIME[5]_net_1 , 
        \timecount_8_iv_2[6] , \S_DUMPTIME[6]_net_1 , 
        \timecount_RNO_6[6]_net_1 , \timecount_8_iv_1[6] , 
        \PLUSECYCLE[6]_net_1 , \timecount_RNO_5[6]_net_1 , 
        \timecount_8_iv_0[6] , \M_DUMPTIME[6]_net_1 , 
        \timecount_8_iv_2[1] , \S_DUMPTIME[1]_net_1 , \CUTTIME_m[1] , 
        \timecount_8_iv_1[1] , \PLUSECYCLE[1]_net_1 , \PLUSETIME_m[1] , 
        \timecount_8_iv_0[1] , \M_DUMPTIME[1]_net_1 , 
        \timecount_8_iv_2[3] , \S_DUMPTIME[3]_net_1 , \CUTTIME_m[3] , 
        \timecount_8_iv_1[3] , \PLUSECYCLE[3]_net_1 , \PLUSETIME_m[3] , 
        \timecount_8_iv_0[3] , \M_DUMPTIME[3]_net_1 , 
        \timecount_8_0_iv_1[11] , \PLUSETIME[11]_net_1 , \CS[5]_net_1 , 
        \S_DUMPTIME_m[11] , \timecount_8_0_iv_0[11] , 
        \M_DUMPTIME[11]_net_1 , \PLUSECYCLE_m[11] , 
        \timecount_8_0_iv_1[12] , \PLUSETIME[12]_net_1 , 
        \S_DUMPTIME_m[12] , \timecount_8_0_iv_0[12] , 
        \M_DUMPTIME[12]_net_1 , \PLUSECYCLE_m[12] , 
        \timecount_8_0_iv_1[13] , \PLUSETIME[13]_net_1 , 
        \S_DUMPTIME_m[13] , \timecount_8_0_iv_0[13] , 
        \M_DUMPTIME[13]_net_1 , \PLUSECYCLE_m[13] , 
        \timecount_8_0_iv_1[15] , \PLUSETIME[15]_net_1 , 
        \S_DUMPTIME_m[15] , \timecount_8_0_iv_0[15] , 
        \M_DUMPTIME[15]_net_1 , \PLUSECYCLE_m[15] , 
        \timecount_8_0_iv_1[0] , \PLUSETIME[0]_net_1 , 
        \S_DUMPTIME_m[0] , \timecount_8_0_iv_0[0] , 
        \M_DUMPTIME[0]_net_1 , \PLUSECYCLE_m[0] , 
        \timecount_8_0_iv_1[7] , \PLUSETIME[7]_net_1 , 
        \S_DUMPTIME_m[7] , \timecount_8_0_iv_0[7] , 
        \M_DUMPTIME[7]_net_1 , \PLUSECYCLE_m[7] , 
        \timecount_8_0_iv_1[8] , \PLUSETIME[8]_net_1 , 
        \S_DUMPTIME_m[8] , \timecount_8_0_iv_0[8] , 
        \M_DUMPTIME[8]_net_1 , \PLUSECYCLE_m[8] , 
        \timecount_8_0_iv_1[9] , \PLUSETIME[9]_net_1 , 
        \S_DUMPTIME_m[9] , \timecount_8_0_iv_0[9] , 
        \M_DUMPTIME[9]_net_1 , \PLUSECYCLE_m[9] , 
        \timecount_8_0_iv_1[10] , \PLUSETIME[10]_net_1 , 
        \S_DUMPTIME_m[10] , \timecount_8_0_iv_0[10] , 
        \M_DUMPTIME[10]_net_1 , \PLUSECYCLE_m[10] , 
        \timecount_8_0_iv_1[14] , \PLUSETIME[14]_net_1 , 
        \S_DUMPTIME_m[14] , \timecount_8_0_iv_0[14] , 
        \M_DUMPTIME[14]_net_1 , \PLUSECYCLE_m[14] , 
        \timecount_8_0_iv_1[4] , \PLUSETIME[4]_net_1 , 
        \S_DUMPTIME_m[4] , \timecount_8_0_iv_0[4] , 
        \M_DUMPTIME[4]_net_1 , \PLUSECYCLE_m[4] , \CS_srsts_i_0[9] , 
        \CS[8]_net_1 , \CS_srsts_i_0[8] , \CS_srsts_i_0[7] , 
        \CS_srsts_i_0[5] , \CS_srsts_i_0[2] , \CS[2]_net_1 , 
        N_290s_i_i_0, \CS_srsts_i_0[3] , \CS[3]_net_1 , 
        \CS_srsts_i_0[4] , \CS_srsts_i_0[6] , \CS_srsts_i_0[1] , 
        \CS[1]_net_1 , un1_PLUSECYCLE14_i_a2_0_net_1, \timecount_8[4] , 
        \CUTTIME_m[4] , \timecount_8[14] , \CUTTIME_m[14] , 
        \timecount_8[10] , \CUTTIME_m[10] , \timecount_8[9] , 
        \CUTTIME_m[9] , \timecount_8[8] , \CUTTIME_m[8] , 
        \timecount_8[7] , \CUTTIME_m[7] , \timecount_8_iv_i_0[6] , 
        \timecount_8_iv_i_0[5] , \timecount_8[3] , 
        \timecount_8_iv_i_0[2] , \timecount_8[0] , \CUTTIME_m[0] , 
        N_341, N_342_1, \timecount_8[15] , \CUTTIME_m[15] , 
        \timecount_8[13] , \CUTTIME_m[13] , \timecount_8[12] , 
        \CUTTIME_m[12] , \timecount_8[11] , \CUTTIME_m[11] , 
        \CS_RNO_1[6] , \CS_RNO_1[5] , \CS_RNO_1[4] , \CS_RNO_1[3] , 
        \CS_RNO_0[8]_net_1 , \CS_RNO_1[7] , M_DUMPTIME_1_sqmuxa, N_17, 
        PLUSECYCLE_0_sqmuxa, PLUSETIME_1_sqmuxa, S_DUMPTIME_1_sqmuxa, 
        \CS_i_RNO_0[0]_net_1 , \CS[9]_net_1 , \CS_RNO_1[1] , 
        \CS_RNO_1[2] , \CS_RNO_0[9]_net_1 , \timecount_8[1] , N_89, 
        N_343, N_154, N_342, N_155, N_157, N_340, N_158, N_69, N_71, 
        N_72, N_73, N_74, N_75, N_76, N_77, N_78, N_79, N_80, N_81, 
        N_82, N_83, N_84, N_85, \timecount_8[16] , N_87, 
        \timecount_8[18] , N_88, \timecount_8[19] , N_16, 
        \PLUSECYCLE[4]_net_1 , \S_DUMPTIME[4]_net_1 , 
        \CUTTIME[4]_net_1 , \CUTTIME[16]_net_1 , \CUTTIME[18]_net_1 , 
        \CUTTIME[19]_net_1 , \PLUSECYCLE[0]_net_1 , 
        \S_DUMPTIME[0]_net_1 , \CUTTIME[0]_net_1 , 
        \PLUSETIME[2]_net_1 , \CUTTIME[2]_net_1 , \PLUSETIME[3]_net_1 , 
        \CUTTIME[3]_net_1 , \PLUSETIME[5]_net_1 , \CUTTIME[5]_net_1 , 
        \PLUSETIME[6]_net_1 , \CUTTIME[6]_net_1 , 
        \PLUSECYCLE[7]_net_1 , \S_DUMPTIME[7]_net_1 , 
        \CUTTIME[7]_net_1 , \PLUSECYCLE[8]_net_1 , 
        \S_DUMPTIME[8]_net_1 , \CUTTIME[8]_net_1 , 
        \PLUSECYCLE[9]_net_1 , \S_DUMPTIME[9]_net_1 , 
        \CUTTIME[9]_net_1 , \PLUSECYCLE[10]_net_1 , 
        \S_DUMPTIME[10]_net_1 , \CUTTIME[10]_net_1 , 
        \PLUSECYCLE[14]_net_1 , \S_DUMPTIME[14]_net_1 , 
        \CUTTIME[14]_net_1 , \PLUSECYCLE[11]_net_1 , 
        \S_DUMPTIME[11]_net_1 , \CUTTIME[11]_net_1 , 
        \PLUSECYCLE[12]_net_1 , \S_DUMPTIME[12]_net_1 , 
        \CUTTIME[12]_net_1 , \PLUSECYCLE[13]_net_1 , 
        \S_DUMPTIME[13]_net_1 , \CUTTIME[13]_net_1 , 
        \PLUSECYCLE[15]_net_1 , \S_DUMPTIME[15]_net_1 , 
        \CUTTIME[15]_net_1 , bri_cycle_RNO_0_net_1, 
        pluse_start_RNO_1_net_1, rt_sw_RNO_1, soft_dump_RNO_net_1, 
        dump_start_RNO_1_net_1, \timecount_RNO[2]_net_1 , 
        \timecount_RNO[3]_net_1 , \timecount_RNO[4]_net_1 , 
        \timecount_RNO[5]_net_1 , \timecount_RNO[6]_net_1 , 
        \timecount_RNO[7]_net_1 , \timecount_RNO[8]_net_1 , 
        \timecount_RNO[9]_net_1 , \timecount_RNO[10]_net_1 , 
        \timecount_RNO[11]_net_1 , \timecount_RNO[12]_net_1 , 
        \timecount_RNO[13]_net_1 , \timecount_RNO[14]_net_1 , 
        \timecount_RNO[15]_net_1 , \timecount_RNO[16]_net_1 , 
        \timecount_RNO[18]_net_1 , \timecount_RNO[19]_net_1 , 
        \timecount_RNO[0]_net_1 , N_366_i, N_398, 
        \timecount_RNO[17]_net_1 , N_86, \timecount_RNO[1]_net_1 , 
        N_70, reset_out_RNO_0_net_1, N_156, \CUTTIME[1]_net_1 , 
        \PLUSETIME[1]_net_1 , \timecount_8[17] , \CUTTIME[17]_net_1 , 
        GND, VCC, GND_0, VCC_0;
    
    MX2 \timecount_RNO_0[16]  (.A(\timecount_8[16] ), .B(
        timecount_0[16]), .S(\CS[9]_net_1 ), .Y(N_85));
    NOR2B dump_start_RNO (.A(top_code_0_state_1ms_rst_n_0), .B(N_89), 
        .Y(dump_start_RNO_1_net_1));
    OR3C \timecount_RNO_1[4]  (.A(\timecount_8_0_iv_0[4] ), .B(
        \CUTTIME_m[4] ), .C(\timecount_8_0_iv_1[4] ), .Y(
        \timecount_8[4] ));
    DFN1E0 \CUTTIME[2]  (.D(state_1ms_data[2]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[2]_net_1 ));
    MX2 \timecount_RNO_0[1]  (.A(\timecount_8[1] ), .B(timecount_0[1]), 
        .S(\CS[9]_net_1 ), .Y(N_70));
    DFN1E1 \M_DUMPTIME[4]  (.D(state_1ms_data[4]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[4]_net_1 ));
    DFN1E1 \PLUSETIME[12]  (.D(state_1ms_data[12]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[12]_net_1 ));
    DFN1 \timecount[13]  (.D(\timecount_RNO[13]_net_1 ), .CLK(GLA), .Q(
        timecount_0[13]));
    DFN1 \timecount[14]  (.D(\timecount_RNO[14]_net_1 ), .CLK(GLA), .Q(
        timecount_0[14]));
    DFN1E0 \CUTTIME[9]  (.D(state_1ms_data[9]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[9]_net_1 ));
    AOI1B \timecount_RNO_4[9]  (.A(\PLUSETIME[9]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[9] ), .Y(
        \timecount_8_0_iv_1[9] ));
    DFN1E1 \S_DUMPTIME[0]  (.D(state_1ms_data[0]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[0]_net_1 ));
    DFN1E0 \CUTTIME[0]  (.D(state_1ms_data[0]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[0]_net_1 ));
    DFN1E1 \S_DUMPTIME[6]  (.D(state_1ms_data[6]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[6]_net_1 ));
    DFN1E1 \PLUSETIME[11]  (.D(state_1ms_data[11]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[11]_net_1 ));
    OR2B \timecount_RNO_3[0]  (.A(\CUTTIME[0]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[0] ));
    DFN1E1 \PLUSETIME[9]  (.D(state_1ms_data[9]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[9]_net_1 ));
    DFN1E1 \M_DUMPTIME[11]  (.D(state_1ms_data[11]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[11]_net_1 ));
    DFN1E0 \CUTTIME[6]  (.D(state_1ms_data[6]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[6]_net_1 ));
    OA1C \CS_RNO[4]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[3]_net_1 ), 
        .C(\CS_srsts_i_0[4] ), .Y(\CS_RNO_1[4] ));
    NOR2B reset_out_RNO (.A(top_code_0_state_1ms_rst_n), .B(N_156), .Y(
        reset_out_RNO_0_net_1));
    NOR2B rt_sw_RNO (.A(top_code_0_state_1ms_rst_n_0), .B(N_155), .Y(
        rt_sw_RNO_1));
    OR2A \timecount_RNO[0]  (.A(top_code_0_state_1ms_rst_n), .B(N_69), 
        .Y(\timecount_RNO[0]_net_1 ));
    OR2 \CS_RNI5A99[1]  (.A(\CS[8]_net_1 ), .B(\CS[1]_net_1 ), .Y(
        N_342_1));
    DFN1E0 \CUTTIME[16]  (.D(state_1ms_data[0]), .CLK(GLA), .E(N_398), 
        .Q(\CUTTIME[16]_net_1 ));
    OA1B \CS_RNO[9]  (.A(\CS[9]_net_1 ), .B(timer_top_0_clk_en_st1ms), 
        .C(\CS_srsts_i_0[9] ), .Y(\CS_RNO_0[9]_net_1 ));
    DFN1E1 \S_DUMPTIME[1]  (.D(state_1ms_data[1]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[1]_net_1 ));
    MX2 \timecount_RNO_0[8]  (.A(\timecount_8[8] ), .B(timecount_0[8]), 
        .S(\CS[9]_net_1 ), .Y(N_77));
    OA1A \timecount_RNO_4[2]  (.A(\CS[7]_net_1 ), .B(
        \S_DUMPTIME[2]_net_1 ), .C(\timecount_RNO_6[2]_net_1 ), .Y(
        \timecount_8_iv_2[2] ));
    NOR2 soft_dump_RNO_1 (.A(N_342_1), .B(\CS[2]_net_1 ), .Y(N_342));
    NOR2B \timecount_RNO_1[18]  (.A(\CUTTIME[18]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\timecount_8[18] ));
    MX2 \timecount_RNO_0[6]  (.A(\timecount_8_iv_i_0[6] ), .B(
        timecount_0[6]), .S(\CS[9]_net_1 ), .Y(N_75));
    DFN1 \CS[4]  (.D(\CS_RNO_1[4] ), .CLK(GLA), .Q(\CS[4]_net_1 ));
    NOR2B bri_cycle_RNO (.A(top_code_0_state_1ms_rst_n_0), .B(N_158), 
        .Y(bri_cycle_RNO_0_net_1));
    OR2B \timecount_RNO_6[0]  (.A(\S_DUMPTIME[0]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[0] ));
    DFN1 \timecount[8]  (.D(\timecount_RNO[8]_net_1 ), .CLK(GLA), .Q(
        timecount_0[8]));
    OAI1 \CS_RNO_0[4]  (.A(\CS[4]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[4] ));
    OR2B \timecount_RNO_6[12]  (.A(\S_DUMPTIME[12]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[12] ));
    OR2B \timecount_RNO_5[11]  (.A(\PLUSECYCLE[11]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[11] ));
    AOI1B \timecount_RNO_2[13]  (.A(\M_DUMPTIME[13]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[13] ), .Y(
        \timecount_8_0_iv_0[13] ));
    DFN1 \timecount[11]  (.D(\timecount_RNO[11]_net_1 ), .CLK(GLA), .Q(
        timecount_0[11]));
    DFN1E1 \M_DUMPTIME[10]  (.D(state_1ms_data[10]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[10]_net_1 ));
    OR2B \timecount_RNO_6[1]  (.A(\CUTTIME[1]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[1] ));
    DFN1E0 \CUTTIME[19]  (.D(state_1ms_data[3]), .CLK(GLA), .E(N_398), 
        .Q(\CUTTIME[19]_net_1 ));
    DFN1E1 \S_DUMPTIME[14]  (.D(state_1ms_data[14]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[14]_net_1 ));
    DFN1E1 \PLUSETIME[14]  (.D(state_1ms_data[14]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[14]_net_1 ));
    OR3C \timecount_RNO_1[11]  (.A(\timecount_8_0_iv_0[11] ), .B(
        \CUTTIME_m[11] ), .C(\timecount_8_0_iv_1[11] ), .Y(
        \timecount_8[11] ));
    AOI1B \timecount_RNO_2[10]  (.A(\M_DUMPTIME[10]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[10] ), .Y(
        \timecount_8_0_iv_0[10] ));
    AOI1B \timecount_RNO_2[15]  (.A(\M_DUMPTIME[15]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[15] ), .Y(
        \timecount_8_0_iv_0[15] ));
    DFN1E1 \PLUSETIME[5]  (.D(state_1ms_data[5]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[5]_net_1 ));
    OR2B \timecount_RNO_3[9]  (.A(\CUTTIME[9]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[9] ));
    OR2B \timecount_RNO_5[7]  (.A(\PLUSECYCLE[7]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[7] ));
    DFN1E1 \S_DUMPTIME[8]  (.D(state_1ms_data[8]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[8]_net_1 ));
    DFN1 \CS[3]  (.D(\CS_RNO_1[3] ), .CLK(GLA), .Q(\CS[3]_net_1 ));
    DFN1E1 \PLUSECYCLE[11]  (.D(state_1ms_data[11]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[11]_net_1 ));
    DFN1E0 \CUTTIME[8]  (.D(state_1ms_data[8]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[8]_net_1 ));
    AOI1B \timecount_RNO_4[8]  (.A(\PLUSETIME[8]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[8] ), .Y(
        \timecount_8_0_iv_1[8] ));
    AOI1B \timecount_RNO_3[1]  (.A(\M_DUMPTIME[1]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\CS_i[0]_net_1 ), .Y(\timecount_8_iv_0[1] ));
    OA1C \CS_RNO[5]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[4]_net_1 ), 
        .C(\CS_srsts_i_0[5] ), .Y(\CS_RNO_1[5] ));
    DFN1 \timecount[2]  (.D(\timecount_RNO[2]_net_1 ), .CLK(GLA), .Q(
        timecount_0[2]));
    OAI1 \CS_RNO_0[5]  (.A(\CS[5]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[5] ));
    OR2B \timecount_RNO_6[14]  (.A(\S_DUMPTIME[14]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[14] ));
    OA1A \timecount_RNO_2[6]  (.A(\CS[4]_net_1 ), .B(
        \PLUSECYCLE[6]_net_1 ), .C(\timecount_RNO_5[6]_net_1 ), .Y(
        \timecount_8_iv_1[6] ));
    MX2 \timecount_RNO_0[3]  (.A(\timecount_8[3] ), .B(timecount_0[3]), 
        .S(\CS[9]_net_1 ), .Y(N_72));
    DFN1E1 \PLUSETIME[15]  (.D(state_1ms_data[15]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[15]_net_1 ));
    DFN1E1 \M_DUMPTIME[12]  (.D(state_1ms_data[12]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[12]_net_1 ));
    MX2A \CS_RNO_0[1]  (.A(\CS[1]_net_1 ), .B(\CS_i[0]_net_1 ), .S(
        timer_top_0_clk_en_st1ms), .Y(\CS_srsts_i_0[1] ));
    NOR3C S_DUMPTIME_1_sqmuxa_0_a2 (.A(state_1ms_lc[0]), .B(
        state_1ms_lc[1]), .C(N_17), .Y(S_DUMPTIME_1_sqmuxa));
    AOI1B \timecount_RNO_4[13]  (.A(\PLUSETIME[13]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[13] ), .Y(
        \timecount_8_0_iv_1[13] ));
    OR2B \timecount_RNO_3[7]  (.A(\CUTTIME[7]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[7] ));
    OR2B \timecount_RNO_3[11]  (.A(\CUTTIME[11]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[11] ));
    DFN1E1 \PLUSETIME[8]  (.D(state_1ms_data[8]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[8]_net_1 ));
    AOI1B \timecount_RNO_4[4]  (.A(\PLUSETIME[4]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[4] ), .Y(
        \timecount_8_0_iv_1[4] ));
    DFN1 \CS[1]  (.D(\CS_RNO_1[1] ), .CLK(GLA), .Q(\CS[1]_net_1 ));
    NOR3A PLUSECYCLE_0_sqmuxa_0_a2 (.A(N_17), .B(state_1ms_lc[0]), .C(
        state_1ms_lc[1]), .Y(PLUSECYCLE_0_sqmuxa));
    AOI1B \timecount_RNO_2[0]  (.A(\M_DUMPTIME[0]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[0] ), .Y(
        \timecount_8_0_iv_0[0] ));
    NOR2B \timecount_RNO[12]  (.A(top_code_0_state_1ms_rst_n), .B(N_81)
        , .Y(\timecount_RNO[12]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1 \PLUSETIME[10]  (.D(state_1ms_data[10]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[10]_net_1 ));
    NOR2B \timecount_RNO[9]  (.A(top_code_0_state_1ms_rst_n), .B(N_78), 
        .Y(\timecount_RNO[9]_net_1 ));
    DFN1E1 \PLUSECYCLE[7]  (.D(state_1ms_data[7]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[7]_net_1 ));
    DFN1E0 \CUTTIME[3]  (.D(state_1ms_data[3]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[3]_net_1 ));
    DFN1 bri_cycle (.D(bri_cycle_RNO_0_net_1), .CLK(GLA), .Q(
        state_1ms_0_bri_cycle));
    AOI1 \CS_i_RNO[0]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[9]_net_1 )
        , .C(N_290s_i_i_0), .Y(\CS_i_RNO_0[0]_net_1 ));
    MX2 dump_start_RNO_0 (.A(state_1ms_0_dump_start), .B(N_341), .S(
        N_343), .Y(N_89));
    DFN1 \CS_i[0]  (.D(\CS_i_RNO_0[0]_net_1 ), .CLK(GLA), .Q(
        \CS_i[0]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    AOI1B \timecount_RNO_4[10]  (.A(\PLUSETIME[10]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[10] ), .Y(
        \timecount_8_0_iv_1[10] ));
    AOI1B \timecount_RNO_4[15]  (.A(\PLUSETIME[15]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[15] ), .Y(
        \timecount_8_0_iv_1[15] ));
    MX2 \timecount_RNO_0[13]  (.A(\timecount_8[13] ), .B(
        timecount_0[13]), .S(\CS[9]_net_1 ), .Y(N_82));
    NOR3B PLUSETIME_1_sqmuxa_0_a2 (.A(state_1ms_lc[0]), .B(N_17), .C(
        state_1ms_lc[1]), .Y(PLUSETIME_1_sqmuxa));
    MX2 soft_dump_RNO_0 (.A(state_1ms_0_soft_dump), .B(N_342), .S(
        N_343), .Y(N_154));
    OA1C \CS_RNO[7]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[6]_net_1 ), 
        .C(\CS_srsts_i_0[7] ), .Y(\CS_RNO_1[7] ));
    DFN1 \timecount[9]  (.D(\timecount_RNO[9]_net_1 ), .CLK(GLA), .Q(
        timecount_0[9]));
    OR3C \timecount_RNO_1[3]  (.A(\timecount_8_iv_1[3] ), .B(
        \timecount_8_iv_0[3] ), .C(\timecount_8_iv_2[3] ), .Y(
        \timecount_8[3] ));
    OR2B \timecount_RNO_5[12]  (.A(\PLUSECYCLE[12]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[12] ));
    DFN1E0 \CUTTIME[15]  (.D(state_1ms_data[15]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[15]_net_1 ));
    DFN1E1 \PLUSECYCLE[14]  (.D(state_1ms_data[14]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[14]_net_1 ));
    MX2 \timecount_RNO_0[10]  (.A(\timecount_8[10] ), .B(
        timecount_0[10]), .S(\CS[9]_net_1 ), .Y(N_79));
    MX2 \timecount_RNO_0[15]  (.A(\timecount_8[15] ), .B(
        timecount_0[15]), .S(\CS[9]_net_1 ), .Y(N_84));
    DFN1E1 \M_DUMPTIME[7]  (.D(state_1ms_data[7]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[7]_net_1 ));
    MX2 \timecount_RNO_0[19]  (.A(\timecount_8[19] ), .B(
        timecount_0[19]), .S(\CS[9]_net_1 ), .Y(N_88));
    DFN1E1 \PLUSETIME[3]  (.D(state_1ms_data[3]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[3]_net_1 ));
    OR3C \timecount_RNO_1[12]  (.A(\timecount_8_0_iv_0[12] ), .B(
        \CUTTIME_m[12] ), .C(\timecount_8_0_iv_1[12] ), .Y(
        \timecount_8[12] ));
    DFN1 \timecount[12]  (.D(\timecount_RNO[12]_net_1 ), .CLK(GLA), .Q(
        timecount_0[12]));
    OR2B \timecount_RNO_6[7]  (.A(\S_DUMPTIME[7]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[7] ));
    OA1C \CS_RNO[3]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[2]_net_1 ), 
        .C(\CS_srsts_i_0[3] ), .Y(\CS_RNO_1[3] ));
    MX2 \timecount_RNO_0[9]  (.A(\timecount_8[9] ), .B(timecount_0[9]), 
        .S(\CS[9]_net_1 ), .Y(N_78));
    DFN1E1 \PLUSETIME[4]  (.D(state_1ms_data[4]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[4]_net_1 ));
    DFN1 \timecount[7]  (.D(\timecount_RNO[7]_net_1 ), .CLK(GLA), .Q(
        timecount_0[7]));
    OR2B \timecount_RNO_5[3]  (.A(\PLUSETIME[3]_net_1 ), .B(
        \CS[5]_net_1 ), .Y(\PLUSETIME_m[3] ));
    MX2B reset_out_RNO_0 (.A(state_1ms_0_reset_out), .B(\CS[1]_net_1 ), 
        .S(N_343), .Y(N_156));
    DFN1E1 \PLUSECYCLE[5]  (.D(state_1ms_data[5]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[5]_net_1 ));
    OAI1 \CS_RNO_0[6]  (.A(\CS[6]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[6] ));
    NOR2A \CS_RNO[1]  (.A(top_code_0_state_1ms_rst_n_0), .B(
        \CS_srsts_i_0[1] ), .Y(\CS_RNO_1[1] ));
    DFN1E1 \M_DUMPTIME[3]  (.D(state_1ms_data[3]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[3]_net_1 ));
    DFN1 \timecount[19]  (.D(\timecount_RNO[19]_net_1 ), .CLK(GLA), .Q(
        timecount_0[19]));
    DFN1 \CS[9]  (.D(\CS_RNO_0[9]_net_1 ), .CLK(GLA), .Q(\CS[9]_net_1 )
        );
    VCC VCC_i (.Y(VCC));
    DFN1E1 \S_DUMPTIME[2]  (.D(state_1ms_data[2]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[2]_net_1 ));
    MX2 \timecount_RNO_0[4]  (.A(\timecount_8[4] ), .B(timecount_0[4]), 
        .S(\CS[9]_net_1 ), .Y(N_73));
    OR2A un1_PLUSECYCLE14_i_a2_0 (.A(top_code_0_state_1ms_load), .B(
        state_1ms_lc[3]), .Y(N_16));
    OR2A \timecount_RNO_6[6]  (.A(\CS[8]_net_1 ), .B(
        \CUTTIME[6]_net_1 ), .Y(\timecount_RNO_6[6]_net_1 ));
    DFN1E1 \S_DUMPTIME[5]  (.D(state_1ms_data[5]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[5]_net_1 ));
    DFN1E0 \CUTTIME[11]  (.D(state_1ms_data[11]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[11]_net_1 ));
    OR2B \timecount_RNO_5[14]  (.A(\PLUSECYCLE[14]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[14] ));
    DFN1E1 \M_DUMPTIME[14]  (.D(state_1ms_data[14]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[14]_net_1 ));
    OA1A \timecount_RNO_3[2]  (.A(\CS[6]_net_1 ), .B(
        \M_DUMPTIME[2]_net_1 ), .C(\CS_i[0]_net_1 ), .Y(
        \timecount_8_iv_0[2] ));
    OAI1 \CS_RNO_0[2]  (.A(\CS[2]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[2] ));
    MX2 bri_cycle_RNO_0 (.A(state_1ms_0_bri_cycle), .B(\CS[5]_net_1 ), 
        .S(N_343), .Y(N_158));
    DFN1E1 \PLUSECYCLE[4]  (.D(state_1ms_data[4]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[4]_net_1 ));
    NOR2B \timecount_RNO[16]  (.A(top_code_0_state_1ms_rst_n), .B(N_85)
        , .Y(\timecount_RNO[16]_net_1 ));
    OR2B \timecount_RNO_3[12]  (.A(\CUTTIME[12]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[12] ));
    MX2 rt_sw_RNO_0 (.A(state_1ms_0_rt_sw), .B(\CS[7]_net_1 ), .S(
        N_343), .Y(N_155));
    DFN1 \timecount[6]  (.D(\timecount_RNO[6]_net_1 ), .CLK(GLA), .Q(
        timecount_0[6]));
    OR3C \timecount_RNO_1[9]  (.A(\timecount_8_0_iv_0[9] ), .B(
        \CUTTIME_m[9] ), .C(\timecount_8_0_iv_1[9] ), .Y(
        \timecount_8[9] ));
    DFN1E1 \PLUSECYCLE[8]  (.D(state_1ms_data[8]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[8]_net_1 ));
    OR2B \timecount_RNO_6[9]  (.A(\S_DUMPTIME[9]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[9] ));
    OR3C \timecount_RNO_1[14]  (.A(\timecount_8_0_iv_0[14] ), .B(
        \CUTTIME_m[14] ), .C(\timecount_8_0_iv_1[14] ), .Y(
        \timecount_8[14] ));
    MX2 \timecount_RNO_0[0]  (.A(\timecount_8[0] ), .B(timecount_0[0]), 
        .S(\CS[9]_net_1 ), .Y(N_69));
    NOR2B pluse_start_RNO (.A(top_code_0_state_1ms_rst_n_0), .B(N_157), 
        .Y(pluse_start_RNO_1_net_1));
    NOR2B \timecount_RNO[17]  (.A(top_code_0_state_1ms_rst_n), .B(N_86)
        , .Y(\timecount_RNO[17]_net_1 ));
    MX2 \timecount_RNO_0[17]  (.A(\timecount_8[17] ), .B(
        timecount_0[17]), .S(\CS[9]_net_1 ), .Y(N_86));
    DFN1 \timecount[15]  (.D(\timecount_RNO[15]_net_1 ), .CLK(GLA), .Q(
        timecount_0[15]));
    NOR2 S_DUMPTIME_1_sqmuxa_0_a2_0 (.A(state_1ms_lc[2]), .B(N_16), .Y(
        N_17));
    NOR2B \timecount_RNO[5]  (.A(top_code_0_state_1ms_rst_n_0), .B(
        N_74), .Y(\timecount_RNO[5]_net_1 ));
    OR2B \timecount_RNO_6[4]  (.A(\S_DUMPTIME[4]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[4] ));
    DFN1E1 \PLUSECYCLE[2]  (.D(state_1ms_data[2]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[2]_net_1 ));
    OA1A \timecount_RNO_4[6]  (.A(\CS[7]_net_1 ), .B(
        \S_DUMPTIME[6]_net_1 ), .C(\timecount_RNO_6[6]_net_1 ), .Y(
        \timecount_8_iv_2[6] ));
    NOR3 dump_start_RNO_1 (.A(\CS[7]_net_1 ), .B(\CS[2]_net_1 ), .C(
        N_342_1), .Y(N_341));
    NOR3C \timecount_RNO_1[6]  (.A(\timecount_8_iv_1[6] ), .B(
        \timecount_8_iv_0[6] ), .C(\timecount_8_iv_2[6] ), .Y(
        \timecount_8_iv_i_0[6] ));
    DFN1E1 \M_DUMPTIME[15]  (.D(state_1ms_data[15]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[15]_net_1 ));
    DFN1E1 \M_DUMPTIME[0]  (.D(state_1ms_data[0]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[0]_net_1 ));
    OR2B \timecount_RNO_5[1]  (.A(\PLUSETIME[1]_net_1 ), .B(
        \CS[5]_net_1 ), .Y(\PLUSETIME_m[1] ));
    DFN1 \timecount[1]  (.D(\timecount_RNO[1]_net_1 ), .CLK(GLA), .Q(
        timecount_0[1]));
    DFN1E1 \M_DUMPTIME[6]  (.D(state_1ms_data[6]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[6]_net_1 ));
    OR2A \timecount_RNO_5[6]  (.A(\CS[5]_net_1 ), .B(
        \PLUSETIME[6]_net_1 ), .Y(\timecount_RNO_5[6]_net_1 ));
    OR2B \timecount_RNO_3[14]  (.A(\CUTTIME[14]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[14] ));
    DFN1 \timecount[10]  (.D(\timecount_RNO[10]_net_1 ), .CLK(GLA), .Q(
        timecount_0[10]));
    AOI1B \timecount_RNO_2[11]  (.A(\M_DUMPTIME[11]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[11] ), .Y(
        \timecount_8_0_iv_0[11] ));
    AO1C \CS_RNO_0[9]  (.A(\CS[8]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[9] ));
    NOR2B \timecount_RNO[3]  (.A(top_code_0_state_1ms_rst_n_0), .B(
        N_72), .Y(\timecount_RNO[3]_net_1 ));
    NOR2B \timecount_RNO[19]  (.A(top_code_0_state_1ms_rst_n), .B(N_88)
        , .Y(\timecount_RNO[19]_net_1 ));
    DFN1 \timecount[18]  (.D(\timecount_RNO[18]_net_1 ), .CLK(GLA), .Q(
        timecount_0[18]));
    NOR2B \timecount_RNO[14]  (.A(top_code_0_state_1ms_rst_n), .B(N_83)
        , .Y(\timecount_RNO[14]_net_1 ));
    DFN1E1 \PLUSECYCLE[1]  (.D(state_1ms_data[1]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[1]_net_1 ));
    DFN1E0 \CUTTIME[5]  (.D(state_1ms_data[5]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[5]_net_1 ));
    DFN1E1 \M_DUMPTIME[1]  (.D(state_1ms_data[1]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[1]_net_1 ));
    NOR3C \timecount_RNO_1[5]  (.A(\timecount_8_iv_1[5] ), .B(
        \timecount_8_iv_0[5] ), .C(\timecount_8_iv_2[5] ), .Y(
        \timecount_8_iv_i_0[5] ));
    DFN1 \timecount[17]  (.D(\timecount_RNO[17]_net_1 ), .CLK(GLA), .Q(
        timecount_0[17]));
    DFN1E1 \PLUSECYCLE[10]  (.D(state_1ms_data[10]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[10]_net_1 ));
    NOR2B \timecount_RNO_1[16]  (.A(\CUTTIME[16]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\timecount_8[16] ));
    MX2 \timecount_RNO_0[5]  (.A(\timecount_8_iv_i_0[5] ), .B(
        timecount_0[5]), .S(\CS[9]_net_1 ), .Y(N_74));
    OA1A \timecount_RNO_4[5]  (.A(\CS[7]_net_1 ), .B(
        \S_DUMPTIME[5]_net_1 ), .C(\timecount_RNO_6[5]_net_1 ), .Y(
        \timecount_8_iv_2[5] ));
    DFN1E1 \S_DUMPTIME[9]  (.D(state_1ms_data[9]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[9]_net_1 ));
    DFN1E0 \CUTTIME[13]  (.D(state_1ms_data[13]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[13]_net_1 ));
    NOR2B \timecount_RNO[13]  (.A(top_code_0_state_1ms_rst_n), .B(N_82)
        , .Y(\timecount_RNO[13]_net_1 ));
    NOR2B \timecount_RNO[1]  (.A(top_code_0_state_1ms_rst_n), .B(N_70), 
        .Y(\timecount_RNO[1]_net_1 ));
    DFN1E1 \S_DUMPTIME[10]  (.D(state_1ms_data[10]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[10]_net_1 ));
    OR2B \timecount_RNO_6[8]  (.A(\S_DUMPTIME[8]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[8] ));
    MX2 \timecount_RNO_0[18]  (.A(\timecount_8[18] ), .B(
        timecount_0[18]), .S(\CS[9]_net_1 ), .Y(N_87));
    DFN1E0 \CUTTIME[17]  (.D(state_1ms_data[1]), .CLK(GLA), .E(N_398), 
        .Q(\CUTTIME[17]_net_1 ));
    NOR2B soft_dump_RNO (.A(top_code_0_state_1ms_rst_n_0), .B(N_154), 
        .Y(soft_dump_RNO_net_1));
    DFN1 \CS[7]  (.D(\CS_RNO_1[7] ), .CLK(GLA), .Q(\CS[7]_net_1 ));
    DFN1E1 \S_DUMPTIME[4]  (.D(state_1ms_data[4]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[4]_net_1 ));
    AOI1B \timecount_RNO_4[11]  (.A(\PLUSETIME[11]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[11] ), .Y(
        \timecount_8_0_iv_1[11] ));
    DFN1 \CS[6]  (.D(\CS_RNO_1[6] ), .CLK(GLA), .Q(\CS[6]_net_1 ));
    AOI1B \timecount_RNO_4[3]  (.A(\S_DUMPTIME[3]_net_1 ), .B(
        \CS[7]_net_1 ), .C(\CUTTIME_m[3] ), .Y(\timecount_8_iv_2[3] ));
    OR2B \timecount_RNO_6[13]  (.A(\S_DUMPTIME[13]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[13] ));
    DFN1E1 \S_DUMPTIME[15]  (.D(state_1ms_data[15]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[15]_net_1 ));
    AOI1B \timecount_RNO_2[7]  (.A(\M_DUMPTIME[7]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[7] ), .Y(
        \timecount_8_0_iv_0[7] ));
    DFN1E1 \M_DUMPTIME[8]  (.D(state_1ms_data[8]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[8]_net_1 ));
    AOI1B \timecount_RNO_2[8]  (.A(\M_DUMPTIME[8]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[8] ), .Y(
        \timecount_8_0_iv_0[8] ));
    DFN1E0 \CUTTIME[12]  (.D(state_1ms_data[12]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[12]_net_1 ));
    OR3A CUTTIME_81_e (.A(state_1ms_lc[0]), .B(N_16), .C(
        un1_PLUSECYCLE14_i_a2_0_net_1), .Y(N_398));
    MX2 \timecount_RNO_0[11]  (.A(\timecount_8[11] ), .B(
        timecount_0[11]), .S(\CS[9]_net_1 ), .Y(N_80));
    DFN1E0 \CUTTIME[14]  (.D(state_1ms_data[14]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[14]_net_1 ));
    AOI1B \timecount_RNO_2[3]  (.A(\PLUSECYCLE[3]_net_1 ), .B(
        \CS[4]_net_1 ), .C(\PLUSETIME_m[3] ), .Y(\timecount_8_iv_1[3] )
        );
    OR3C \timecount_RNO_1[1]  (.A(\timecount_8_iv_1[1] ), .B(
        \timecount_8_iv_0[1] ), .C(\timecount_8_iv_2[1] ), .Y(
        \timecount_8[1] ));
    OR2B \timecount_RNO_6[10]  (.A(\S_DUMPTIME[10]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[10] ));
    OR2B \timecount_RNO_6[15]  (.A(\S_DUMPTIME[15]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[15] ));
    DFN1 \timecount[16]  (.D(\timecount_RNO[16]_net_1 ), .CLK(GLA), .Q(
        timecount_0[16]));
    DFN1E1 \PLUSECYCLE[9]  (.D(state_1ms_data[9]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[9]_net_1 ));
    OR2B \timecount_RNO_6[3]  (.A(\CUTTIME[3]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[3] ));
    OR2B \timecount_RNO_5[9]  (.A(\PLUSECYCLE[9]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[9] ));
    OR2 pluse_start_RNO_1 (.A(\CS[5]_net_1 ), .B(\CS[4]_net_1 ), .Y(
        N_340));
    OA1C \CS_RNO[2]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[1]_net_1 ), 
        .C(\CS_srsts_i_0[2] ), .Y(\CS_RNO_1[2] ));
    AOI1B \timecount_RNO_4[0]  (.A(\PLUSETIME[0]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[0] ), .Y(
        \timecount_8_0_iv_1[0] ));
    GND GND_i_0 (.Y(GND_0));
    AOI1B \timecount_RNO_2[12]  (.A(\M_DUMPTIME[12]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[12] ), .Y(
        \timecount_8_0_iv_0[12] ));
    DFN1 \CS[8]  (.D(\CS_RNO_0[8]_net_1 ), .CLK(GLA), .Q(\CS[8]_net_1 )
        );
    OR2A un1_PLUSECYCLE14_i_a2_0_0 (.A(state_1ms_lc[2]), .B(
        state_1ms_lc[1]), .Y(un1_PLUSECYCLE14_i_a2_0_net_1));
    DFN1E0 \CUTTIME[7]  (.D(state_1ms_data[7]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[7]_net_1 ));
    AOI1B \timecount_RNO_4[7]  (.A(\PLUSETIME[7]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[7] ), .Y(
        \timecount_8_0_iv_1[7] ));
    OR2B \timecount_RNO_3[8]  (.A(\CUTTIME[8]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[8] ));
    DFN1 \timecount[4]  (.D(\timecount_RNO[4]_net_1 ), .CLK(GLA), .Q(
        timecount_0[4]));
    AO1C \CS_RNO_0[8]  (.A(\CS[7]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[8] ));
    OR2A \timecount_RNO_6[2]  (.A(\CS[8]_net_1 ), .B(
        \CUTTIME[2]_net_1 ), .Y(\timecount_RNO_6[2]_net_1 ));
    OR3C \timecount_RNO_1[8]  (.A(\timecount_8_0_iv_0[8] ), .B(
        \CUTTIME_m[8] ), .C(\timecount_8_0_iv_1[8] ), .Y(
        \timecount_8[8] ));
    DFN1E1 \PLUSECYCLE[0]  (.D(state_1ms_data[0]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[0]_net_1 ));
    NOR2B \timecount_RNO[8]  (.A(top_code_0_state_1ms_rst_n), .B(N_77), 
        .Y(\timecount_RNO[8]_net_1 ));
    OAI1 \CS_i_RNO_0[0]  (.A(\CS_i[0]_net_1 ), .B(
        timer_top_0_clk_en_st1ms), .C(top_code_0_state_1ms_rst_n_0), 
        .Y(N_290s_i_i_0));
    AOI1B \timecount_RNO_2[1]  (.A(\PLUSECYCLE[1]_net_1 ), .B(
        \CS[4]_net_1 ), .C(\PLUSETIME_m[1] ), .Y(\timecount_8_iv_1[1] )
        );
    OR3C \timecount_RNO_1[0]  (.A(\timecount_8_0_iv_0[0] ), .B(
        \CUTTIME_m[0] ), .C(\timecount_8_0_iv_1[0] ), .Y(
        \timecount_8[0] ));
    DFN1 \CS[2]  (.D(\CS_RNO_1[2] ), .CLK(GLA), .Q(\CS[2]_net_1 ));
    OR2A \timecount_RNO_6[5]  (.A(\CS[8]_net_1 ), .B(
        \CUTTIME[5]_net_1 ), .Y(\timecount_RNO_6[5]_net_1 ));
    OR2A \timecount_RNO_5[5]  (.A(\CS[5]_net_1 ), .B(
        \PLUSETIME[5]_net_1 ), .Y(\timecount_RNO_5[5]_net_1 ));
    AOI1B \timecount_RNO_2[14]  (.A(\M_DUMPTIME[14]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[14] ), .Y(
        \timecount_8_0_iv_0[14] ));
    OR2B \timecount_RNO_5[0]  (.A(\PLUSECYCLE[0]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[0] ));
    NOR2B \timecount_RNO[4]  (.A(top_code_0_state_1ms_rst_n_0), .B(
        N_73), .Y(\timecount_RNO[4]_net_1 ));
    DFN1E1 \PLUSECYCLE[3]  (.D(state_1ms_data[3]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[3]_net_1 ));
    DFN1E1 \PLUSECYCLE[12]  (.D(state_1ms_data[12]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[12]_net_1 ));
    AOI1B \timecount_RNO_4[12]  (.A(\PLUSETIME[12]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[12] ), .Y(
        \timecount_8_0_iv_1[12] ));
    DFN1E0 \CUTTIME[18]  (.D(state_1ms_data[2]), .CLK(GLA), .E(N_398), 
        .Q(\CUTTIME[18]_net_1 ));
    OR2B \timecount_RNO_5[13]  (.A(\PLUSECYCLE[13]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[13] ));
    DFN1E1 \PLUSETIME[6]  (.D(state_1ms_data[6]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[6]_net_1 ));
    DFN1E1 \PLUSETIME[13]  (.D(state_1ms_data[13]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[13]_net_1 ));
    DFN1 dump_start (.D(dump_start_RNO_1_net_1), .CLK(GLA), .Q(
        state_1ms_0_dump_start));
    MX2 \timecount_RNO_0[2]  (.A(\timecount_8_iv_i_0[2] ), .B(
        timecount_0[2]), .S(\CS[9]_net_1 ), .Y(N_71));
    DFN1E0 \CUTTIME[10]  (.D(state_1ms_data[10]), .CLK(GLA), .E(
        N_366_i), .Q(\CUTTIME[10]_net_1 ));
    OA1A \timecount_RNO_2[5]  (.A(\CS[4]_net_1 ), .B(
        \PLUSECYCLE[5]_net_1 ), .C(\timecount_RNO_5[5]_net_1 ), .Y(
        \timecount_8_iv_1[5] ));
    NOR2A \CS_i_RNIT6K5[0]  (.A(\CS_i[0]_net_1 ), .B(\CS[9]_net_1 ), 
        .Y(N_343));
    MX2 \timecount_RNO_0[12]  (.A(\timecount_8[12] ), .B(
        timecount_0[12]), .S(\CS[9]_net_1 ), .Y(N_81));
    DFN1E1 \M_DUMPTIME[2]  (.D(state_1ms_data[2]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[2]_net_1 ));
    OR3C \timecount_RNO_1[13]  (.A(\timecount_8_0_iv_0[13] ), .B(
        \CUTTIME_m[13] ), .C(\timecount_8_0_iv_1[13] ), .Y(
        \timecount_8[13] ));
    MX2 pluse_start_RNO_0 (.A(state_1ms_0_pluse_start), .B(N_340), .S(
        N_343), .Y(N_157));
    DFN1E1 \PLUSECYCLE[13]  (.D(state_1ms_data[13]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[13]_net_1 ));
    DFN1E1 \M_DUMPTIME[5]  (.D(state_1ms_data[5]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[5]_net_1 ));
    OR2B \timecount_RNO_5[10]  (.A(\PLUSECYCLE[10]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[10] ));
    NOR2B \timecount_RNO[11]  (.A(top_code_0_state_1ms_rst_n), .B(N_80)
        , .Y(\timecount_RNO[11]_net_1 ));
    OR2B \timecount_RNO_5[15]  (.A(\PLUSECYCLE[15]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[15] ));
    DFN1E1 \S_DUMPTIME[12]  (.D(state_1ms_data[12]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[12]_net_1 ));
    DFN1E0 \CUTTIME[1]  (.D(state_1ms_data[1]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[1]_net_1 ));
    DFN1 soft_dump (.D(soft_dump_RNO_net_1), .CLK(GLA), .Q(
        state_1ms_0_soft_dump));
    OA1A \timecount_RNO_3[6]  (.A(\CS[6]_net_1 ), .B(
        \M_DUMPTIME[6]_net_1 ), .C(\CS_i[0]_net_1 ), .Y(
        \timecount_8_iv_0[6] ));
    DFN1 pluse_start (.D(pluse_start_RNO_1_net_1), .CLK(GLA), .Q(
        state_1ms_0_pluse_start));
    NOR2B \timecount_RNO[2]  (.A(top_code_0_state_1ms_rst_n_0), .B(
        N_71), .Y(\timecount_RNO[2]_net_1 ));
    OR3C \timecount_RNO_1[10]  (.A(\timecount_8_0_iv_0[10] ), .B(
        \CUTTIME_m[10] ), .C(\timecount_8_0_iv_1[10] ), .Y(
        \timecount_8[10] ));
    DFN1 \timecount[0]  (.D(\timecount_RNO[0]_net_1 ), .CLK(GLA), .Q(
        timecount_0[0]));
    OR3C \timecount_RNO_1[15]  (.A(\timecount_8_0_iv_0[15] ), .B(
        \CUTTIME_m[15] ), .C(\timecount_8_0_iv_1[15] ), .Y(
        \timecount_8[15] ));
    DFN1E1 \PLUSETIME[0]  (.D(state_1ms_data[0]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[0]_net_1 ));
    AOI1B \timecount_RNO_4[14]  (.A(\PLUSETIME[14]_net_1 ), .B(
        \CS[5]_net_1 ), .C(\S_DUMPTIME_m[14] ), .Y(
        \timecount_8_0_iv_1[14] ));
    NOR2B \timecount_RNO_1[19]  (.A(\CUTTIME[19]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\timecount_8[19] ));
    MX2 \timecount_RNO_0[7]  (.A(\timecount_8[7] ), .B(timecount_0[7]), 
        .S(\CS[9]_net_1 ), .Y(N_76));
    OR2B \timecount_RNO_3[4]  (.A(\CUTTIME[4]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[4] ));
    OA1B \CS_RNO[8]  (.A(\CS[8]_net_1 ), .B(timer_top_0_clk_en_st1ms), 
        .C(\CS_srsts_i_0[8] ), .Y(\CS_RNO_0[8]_net_1 ));
    AOI1B \timecount_RNO_2[4]  (.A(\M_DUMPTIME[4]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[4] ), .Y(
        \timecount_8_0_iv_0[4] ));
    NOR2B \timecount_RNO[15]  (.A(top_code_0_state_1ms_rst_n), .B(N_84)
        , .Y(\timecount_RNO[15]_net_1 ));
    OR2B \timecount_RNO_3[13]  (.A(\CUTTIME[13]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[13] ));
    DFN1 \CS[5]  (.D(\CS_RNO_1[5] ), .CLK(GLA), .Q(\CS[5]_net_1 ));
    OAI1 \CS_RNO_0[3]  (.A(\CS[3]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[3] ));
    OR2B \timecount_RNO_5[4]  (.A(\PLUSECYCLE[4]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[4] ));
    MX2 \timecount_RNO_0[14]  (.A(\timecount_8[14] ), .B(
        timecount_0[14]), .S(\CS[9]_net_1 ), .Y(N_83));
    DFN1E1 \S_DUMPTIME[7]  (.D(state_1ms_data[7]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[7]_net_1 ));
    DFN1E1 \PLUSETIME[2]  (.D(state_1ms_data[2]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[2]_net_1 ));
    DFN1E1 \M_DUMPTIME[13]  (.D(state_1ms_data[13]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[13]_net_1 ));
    OR3 CUTTIME_65_e (.A(N_16), .B(un1_PLUSECYCLE14_i_a2_0_net_1), .C(
        state_1ms_lc[0]), .Y(N_366_i));
    DFN1E1 \PLUSECYCLE[15]  (.D(state_1ms_data[15]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[15]_net_1 ));
    NOR3B M_DUMPTIME_1_sqmuxa_0_a2 (.A(state_1ms_lc[1]), .B(N_17), .C(
        state_1ms_lc[0]), .Y(M_DUMPTIME_1_sqmuxa));
    OR2B \timecount_RNO_3[10]  (.A(\CUTTIME[10]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[10] ));
    NOR2B \timecount_RNO[18]  (.A(top_code_0_state_1ms_rst_n), .B(N_87)
        , .Y(\timecount_RNO[18]_net_1 ));
    OR2B \timecount_RNO_3[15]  (.A(\CUTTIME[15]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\CUTTIME_m[15] ));
    NOR2B \timecount_RNO[6]  (.A(top_code_0_state_1ms_rst_n), .B(N_75), 
        .Y(\timecount_RNO[6]_net_1 ));
    NOR2B \timecount_RNO[7]  (.A(top_code_0_state_1ms_rst_n), .B(N_76), 
        .Y(\timecount_RNO[7]_net_1 ));
    DFN1 rt_sw (.D(rt_sw_RNO_1), .CLK(GLA), .Q(state_1ms_0_rt_sw));
    DFN1E1 \PLUSETIME[7]  (.D(state_1ms_data[7]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[7]_net_1 ));
    OA1C \CS_RNO[6]  (.A(timer_top_0_clk_en_st1ms), .B(\CS[5]_net_1 ), 
        .C(\CS_srsts_i_0[6] ), .Y(\CS_RNO_1[6] ));
    OR2B \timecount_RNO_5[8]  (.A(\PLUSECYCLE[8]_net_1 ), .B(
        \CS[4]_net_1 ), .Y(\PLUSECYCLE_m[8] ));
    DFN1E1 \S_DUMPTIME[11]  (.D(state_1ms_data[11]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[11]_net_1 ));
    AOI1B \timecount_RNO_4[1]  (.A(\S_DUMPTIME[1]_net_1 ), .B(
        \CS[7]_net_1 ), .C(\CUTTIME_m[1] ), .Y(\timecount_8_iv_2[1] ));
    DFN1E1 \S_DUMPTIME[3]  (.D(state_1ms_data[3]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[3]_net_1 ));
    DFN1E1 \PLUSECYCLE[6]  (.D(state_1ms_data[6]), .CLK(GLA), .E(
        PLUSECYCLE_0_sqmuxa), .Q(\PLUSECYCLE[6]_net_1 ));
    OAI1 \CS_RNO_0[7]  (.A(\CS[7]_net_1 ), .B(timer_top_0_clk_en_st1ms)
        , .C(top_code_0_state_1ms_rst_n_0), .Y(\CS_srsts_i_0[7] ));
    NOR2B \timecount_RNO[10]  (.A(top_code_0_state_1ms_rst_n), .B(N_79)
        , .Y(\timecount_RNO[10]_net_1 ));
    DFN1E0 \CUTTIME[4]  (.D(state_1ms_data[4]), .CLK(GLA), .E(N_366_i), 
        .Q(\CUTTIME[4]_net_1 ));
    NOR3C \timecount_RNO_1[2]  (.A(\timecount_8_iv_1[2] ), .B(
        \timecount_8_iv_0[2] ), .C(\timecount_8_iv_2[2] ), .Y(
        \timecount_8_iv_i_0[2] ));
    DFN1E1 \PLUSETIME[1]  (.D(state_1ms_data[1]), .CLK(GLA), .E(
        PLUSETIME_1_sqmuxa), .Q(\PLUSETIME[1]_net_1 ));
    NOR2B \timecount_RNO_1[17]  (.A(\CUTTIME[17]_net_1 ), .B(
        \CS[8]_net_1 ), .Y(\timecount_8[17] ));
    OR2B \timecount_RNO_6[11]  (.A(\S_DUMPTIME[11]_net_1 ), .B(
        \CS[7]_net_1 ), .Y(\S_DUMPTIME_m[11] ));
    AOI1B \timecount_RNO_2[9]  (.A(\M_DUMPTIME[9]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\PLUSECYCLE_m[9] ), .Y(
        \timecount_8_0_iv_0[9] ));
    OR3C \timecount_RNO_1[7]  (.A(\timecount_8_0_iv_0[7] ), .B(
        \CUTTIME_m[7] ), .C(\timecount_8_0_iv_1[7] ), .Y(
        \timecount_8[7] ));
    OA1A \timecount_RNO_3[5]  (.A(\CS[6]_net_1 ), .B(
        \M_DUMPTIME[5]_net_1 ), .C(\CS_i[0]_net_1 ), .Y(
        \timecount_8_iv_0[5] ));
    OR2A \timecount_RNO_5[2]  (.A(\CS[5]_net_1 ), .B(
        \PLUSETIME[2]_net_1 ), .Y(\timecount_RNO_5[2]_net_1 ));
    DFN1E1 \M_DUMPTIME[9]  (.D(state_1ms_data[9]), .CLK(GLA), .E(
        M_DUMPTIME_1_sqmuxa), .Q(\M_DUMPTIME[9]_net_1 ));
    OA1A \timecount_RNO_2[2]  (.A(\CS[4]_net_1 ), .B(
        \PLUSECYCLE[2]_net_1 ), .C(\timecount_RNO_5[2]_net_1 ), .Y(
        \timecount_8_iv_1[2] ));
    DFN1 reset_out (.D(reset_out_RNO_0_net_1), .CLK(GLA), .Q(
        state_1ms_0_reset_out));
    AOI1B \timecount_RNO_3[3]  (.A(\M_DUMPTIME[3]_net_1 ), .B(
        \CS[6]_net_1 ), .C(\CS_i[0]_net_1 ), .Y(\timecount_8_iv_0[3] ));
    DFN1 \timecount[5]  (.D(\timecount_RNO[5]_net_1 ), .CLK(GLA), .Q(
        timecount_0[5]));
    DFN1 \timecount[3]  (.D(\timecount_RNO[3]_net_1 ), .CLK(GLA), .Q(
        timecount_0[3]));
    DFN1E1 \S_DUMPTIME[13]  (.D(state_1ms_data[13]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[13]_net_1 ));
    
endmodule


module sd_sacq_coder(
       i,
       i_3,
       i_0_0_0,
       i_4,
       sd_sacq_data,
       sd_sacq_choice,
       count_4,
       count_1,
       count,
       ddsclkout_c,
       GLA,
       scalestate_0_long_opentime,
       s_acq180_c,
       top_code_0_sd_sacq_load,
       scalestate_0_s_acq,
       net_27
    );
output [10:4] i;
output [3:2] i_3;
input  i_0_0_0;
output [1:0] i_4;
input  [15:0] sd_sacq_data;
input  [3:0] sd_sacq_choice;
input  [4:0] count_4;
input  [7:5] count_1;
input  [21:8] count;
input  ddsclkout_c;
input  GLA;
input  scalestate_0_long_opentime;
input  s_acq180_c;
input  top_code_0_sd_sacq_load;
input  scalestate_0_s_acq;
input  net_27;

    wire \i_0_22[10] , \i_0_20[10] , \i_0_19[10] , \un1_count_2_i[0] , 
        \i_0_12[10] , \i_0_11[10] , \i_0_18[10] , \i_0_8[10] , 
        \i_0_7[10] , \i_0_16[10] , \i_0_4[10] , \i_0_3[10] , 
        \i_0_14[10] , N_368_i_i_0, N_364_i_i_0, \i_0_10[10] , 
        \i_0_5[10] , \i_0_6[10] , \i_0_1[10] , \i_0_2[10] , 
        N_360_i_i_0, \i_0_0[10] , N_316_i_i_0, N_348_i_i_0, 
        N_328_i_i_0, N_340_i_i_0, N_304_i_i_0, N_320_i_i_0, 
        \sd_sacq_data7[13]_net_1 , N_344_i_i_0, 
        \sd_sacq_data7[7]_net_1 , N_324_i_i_0, 
        \sd_sacq_data7[20]_net_1 , N_296_i_i_0, 
        \sd_sacq_data7[14]_net_1 , N_352_i_i_0, 
        \sd_sacq_data7[16]_net_1 , N_312_i_i_0, 
        \sd_sacq_data7[17]_net_1 , N_356_i_i_0, 
        \sd_sacq_data7[21]_net_1 , \i_0_0[9] , 
        \un1_count_5_NE_i_a2_14[0] , \un1_count_5_NE_i_a2_6[0] , 
        \un1_count_5_NE_i_a2_5[0] , N_904, \un1_count_5_NE_i_a2_13[0] , 
        \un1_count_5_NE_i_a2_4[0] , \un1_count_5_NE_i_a2_3[0] , 
        \un1_count_5_NE_i_a2_9[0] , \un1_count_5_NE_i_a2_12[0] , 
        N_404_i_i_0, N_384_i_i_0, \un1_count_5_NE_i_a2_8[0] , 
        N_383_i_i_0, N_409_i_i_0, \un1_count_5_NE_i_a2_2[0] , 
        \sd_sacq_data3[0]_net_1 , \un1_count_5_NE_i_a2_0[0]_net_1 , 
        \sd_sacq_data3[10]_net_1 , N_411_i_i_0, 
        \sd_sacq_data3[1]_net_1 , N_405_i_i_0, 
        \sd_sacq_data3[12]_net_1 , N_382_i_i_0, 
        \sd_sacq_data3[7]_net_1 , N_410_i_i_0, 
        \sd_sacq_data3[13]_net_1 , N_402_i_i_0, 
        \sd_sacq_data3[14]_net_1 , \un1_count_4_NE_i_a2_14[0] , 
        \un1_count_4_NE_i_a2_6[0] , \un1_count_4_NE_i_a2_5[0] , 
        \un1_count_4_NE_i_a2_13[0] , \un1_count_4_NE_i_a2_2[0] , 
        \un1_count_4_NE_i_a2_1[0] , \un1_count_4_NE_i_a2_10[0] , 
        \un1_count_4_NE_i_a2_12[0] , N_394_i_i_0, N_389_i_i_0, 
        \un1_count_4_NE_i_a2_8[0] , N_415_i_i_0, N_393_i_i_0, 
        \un1_count_4_NE_i_a2_4[0] , \sd_sacq_data2[0]_net_1 , 
        \un1_count_4_NE_i_a2_0[0] , \sd_sacq_data2[10]_net_1 , 
        N_416_i_i_0, \sd_sacq_data2[1]_net_1 , N_395_i_i_0, 
        \sd_sacq_data2[12]_net_1 , N_388_i_i_0, 
        \sd_sacq_data2[13]_net_1 , N_392_i_i_0, 
        \sd_sacq_data2[8]_net_1 , N_387_i_i_0, 
        \sd_sacq_data2[14]_net_1 , \i_reg18_NE_i_a2_14[0] , 
        \i_reg18_NE_i_a2_6[0] , \i_reg18_NE_i_a2_5[0] , 
        \i_reg18_NE_i_a2_13[0] , \i_reg18_NE_i_a2_2[0] , 
        \i_reg18_NE_i_a2_1[0] , \i_reg18_NE_i_a2_10[0] , 
        \i_reg18_NE_i_a2_12[0] , N_399_i_i_0, N_379_i_i_0, 
        \i_reg18_NE_i_a2_8[0] , N_420_i_i_0, N_398_i_i_0, 
        \i_reg18_NE_i_a2_4[0] , \sd_sacq_data1[0]_net_1 , 
        \i_reg18_NE_i_a2_0[0] , \sd_sacq_data1[10]_net_1 , N_421_i_i_0, 
        \sd_sacq_data1[1]_net_1 , N_400_i_i_0, 
        \sd_sacq_data1[12]_net_1 , N_377_i_i_0, 
        \sd_sacq_data1[13]_net_1 , N_397_i_i_0, 
        \sd_sacq_data1[8]_net_1 , N_378_i_i_0, 
        \sd_sacq_data1[14]_net_1 , \un1_count_NE_19[0] , 
        \un1_count_NE_11[0] , \un1_count_NE_10[0] , 
        \un1_count_NE_17[0] , \un1_count_NE_18[0] , 
        \un1_count_NE_7[0] , \un1_count_NE_6[0] , \un1_count_NE_15[0] , 
        \un1_count_NE_3[0] , \un1_count_NE_2[0] , \un1_count_NE_13[0] , 
        N_361_i_i, N_337_i_i, \un1_count_NE_9[0] , N_305_i_i, 
        N_293_i_i, \un1_count_NE_5[0] , N_373_i_i, N_297_i_i, 
        \un1_count_NE_1[0] , \sd_sacq_data4[3]_net_1 , N_357_i_i, 
        \sd_sacq_data4[4]_net_1 , N_313_i_i, \sd_sacq_data4[10]_net_1 , 
        N_325_i_i, \sd_sacq_data4[2]_net_1 , N_301_i_i, N_321_i_i, 
        N_329_i_i, N_349_i_i, \un1_count_20_i[0] , N_309_i_i, 
        N_333_i_i, N_353_i_i, N_369_i_i, \un1_count_1_NE_18[0] , 
        \un1_count_1_NE_7[0] , \un1_count_1_NE_6[0] , 
        \un1_count_1_NE_15[0] , \un1_count_1_NE_17[0] , 
        \un1_count_1_NE_3[0] , \un1_count_1_NE_2[0] , 
        \un1_count_1_NE_13[0] , \un1_count_1_NE_16[0] , 
        \un1_count_1_NE_1[0] , \un1_count_1_NE_0[0] , 
        \un1_count_1_NE_10[0] , N_362_i_i, N_338_i_i, 
        \un1_count_1_NE_9[0] , N_306_i_i, N_294_i_i, 
        \un1_count_1_NE_5[0] , \sd_sacq_data5[3]_net_1 , N_358_i_i, 
        \sd_sacq_data5[4]_net_1 , N_314_i_i, \sd_sacq_data5[10]_net_1 , 
        N_326_i_i, \sd_sacq_data5[2]_net_1 , N_302_i_i, 
        \sd_sacq_data5[11]_net_1 , N_330_i_i, 
        \sd_sacq_data5[18]_net_1 , \un1_count_1_20_i[0] , 
        \sd_sacq_data5[8]_net_1 , N_334_i_i, \sd_sacq_data5[19]_net_1 , 
        N_370_i_i, \sd_sacq_data5[21]_net_1 , N_374_i_i, 
        \un1_count_2_NE_18[0] , \un1_count_2_NE_7[0] , 
        \un1_count_2_NE_6[0] , \un1_count_2_NE_15[0] , 
        \un1_count_2_NE_17[0] , \un1_count_2_NE_3[0] , 
        \un1_count_2_NE_2[0] , \un1_count_2_NE_13[0] , 
        \un1_count_2_NE_16[0] , \un1_count_2_NE_1[0] , 
        \un1_count_2_NE_0[0] , \un1_count_2_NE_10[0] , N_363_i_i, 
        N_339_i_i, \un1_count_2_NE_9[0] , N_307_i_i, N_295_i_i, 
        \un1_count_2_NE_5[0] , \sd_sacq_data6[3]_net_1 , N_359_i_i, 
        \sd_sacq_data6[4]_net_1 , N_315_i_i, \sd_sacq_data6[10]_net_1 , 
        N_327_i_i, \sd_sacq_data6[2]_net_1 , N_303_i_i, 
        \sd_sacq_data6[11]_net_1 , N_331_i_i, 
        \sd_sacq_data6[18]_net_1 , \un1_count_2_20_i[0] , 
        \sd_sacq_data6[8]_net_1 , N_335_i_i, \sd_sacq_data6[19]_net_1 , 
        N_371_i_i, \sd_sacq_data6[21]_net_1 , N_375_i_i, 
        \un1_count_5_NE_i_a2_0_2[0]_net_1 , 
        un1_sd_sacq_data117_2_i_a2_0_net_1, 
        un1_sd_sacq_data117_3_i_a2_0_net_1, \i_RNO[5]_net_1 , N_579, 
        N_578_i, \i_RNO[6]_net_1 , N_577, un1_i_reg18_1, 
        \i_RNO[7]_net_1 , un1_count_6, \un1_count_NE[0] , 
        \i_RNO[8]_net_1 , \un1_count_1_NE[0] , un1_count_8, 
        \i_RNO[9]_net_1 , \i_RNO[10]_net_1 , sd_sacq_data1_0_sqmuxa, 
        un1_sd_sacq_data117_1_i_a2_0, N_580, sd_sacq_data2_1_sqmuxa, 
        N_792, sd_sacq_data3_1_sqmuxa, \sd_sacq_data4[20]_net_1 , 
        \sd_sacq_data5[20]_net_1 , \sd_sacq_data6[20]_net_1 , 
        \i_RNO_1[0] , \i_RNO[4]_net_1 , \sd_sacq_data4[5]_net_1 , 
        \sd_sacq_data5[5]_net_1 , \sd_sacq_data6[5]_net_1 , 
        \sd_sacq_data7[5]_net_1 , \sd_sacq_data4[21]_net_1 , 
        \sd_sacq_data4[6]_net_1 , \sd_sacq_data5[6]_net_1 , 
        \sd_sacq_data6[6]_net_1 , \sd_sacq_data7[6]_net_1 , 
        \sd_sacq_data4[7]_net_1 , \sd_sacq_data5[7]_net_1 , 
        \sd_sacq_data6[7]_net_1 , \sd_sacq_data4[8]_net_1 , 
        \sd_sacq_data7[8]_net_1 , \sd_sacq_data4[9]_net_1 , 
        \sd_sacq_data5[9]_net_1 , \sd_sacq_data6[9]_net_1 , 
        \sd_sacq_data7[9]_net_1 , \sd_sacq_data7[10]_net_1 , 
        \sd_sacq_data4[11]_net_1 , \sd_sacq_data7[11]_net_1 , 
        \sd_sacq_data4[12]_net_1 , \sd_sacq_data5[12]_net_1 , 
        \sd_sacq_data6[12]_net_1 , \sd_sacq_data7[12]_net_1 , 
        \sd_sacq_data4[13]_net_1 , \sd_sacq_data5[13]_net_1 , 
        \sd_sacq_data6[13]_net_1 , \sd_sacq_data4[14]_net_1 , 
        \sd_sacq_data5[14]_net_1 , \sd_sacq_data6[14]_net_1 , 
        \sd_sacq_data4[15]_net_1 , \sd_sacq_data5[15]_net_1 , 
        \sd_sacq_data6[15]_net_1 , \sd_sacq_data7[15]_net_1 , 
        \sd_sacq_data7[2]_net_1 , \sd_sacq_data7[3]_net_1 , 
        \sd_sacq_data4[18]_net_1 , \sd_sacq_data7[18]_net_1 , 
        \sd_sacq_data4[19]_net_1 , \sd_sacq_data7[19]_net_1 , 
        \sd_sacq_data4[0]_net_1 , \sd_sacq_data5[0]_net_1 , 
        \sd_sacq_data6[0]_net_1 , \sd_sacq_data7[0]_net_1 , 
        \sd_sacq_data4[1]_net_1 , \sd_sacq_data5[1]_net_1 , 
        \sd_sacq_data6[1]_net_1 , \sd_sacq_data7[1]_net_1 , 
        \sd_sacq_data7[4]_net_1 , \sd_sacq_data4[16]_net_1 , 
        \sd_sacq_data5[16]_net_1 , \sd_sacq_data6[16]_net_1 , 
        \sd_sacq_data4[17]_net_1 , \sd_sacq_data5[17]_net_1 , 
        \sd_sacq_data6[17]_net_1 , \sd_sacq_data1[15]_net_1 , 
        \sd_sacq_data1[5]_net_1 , \sd_sacq_data1[3]_net_1 , 
        \sd_sacq_data3[15]_net_1 , \sd_sacq_data3[5]_net_1 , 
        \sd_sacq_data3[3]_net_1 , \sd_sacq_data2[5]_net_1 , 
        \sd_sacq_data2[15]_net_1 , \sd_sacq_data2[3]_net_1 , 
        \sd_sacq_data2[11]_net_1 , \sd_sacq_data2[7]_net_1 , 
        \sd_sacq_data2[9]_net_1 , \sd_sacq_data2[6]_net_1 , 
        \sd_sacq_data1[11]_net_1 , \sd_sacq_data1[7]_net_1 , 
        \sd_sacq_data1[9]_net_1 , \sd_sacq_data1[6]_net_1 , 
        \sd_sacq_data3[11]_net_1 , \sd_sacq_data3[9]_net_1 , 
        \sd_sacq_data3[6]_net_1 , \sd_sacq_data3[8]_net_1 , 
        \sd_sacq_data3[2]_net_1 , \sd_sacq_data3[4]_net_1 , 
        \sd_sacq_data2[2]_net_1 , \sd_sacq_data2[4]_net_1 , 
        \sd_sacq_data1[2]_net_1 , \sd_sacq_data1[4]_net_1 , N_581_i, 
        N_613, N_625_i, N_657, N_683_i, N_573_1, N_701_i, N_713_i, 
        N_745_i, \i_RNO_1[2] , \i_RNO_1[3] , GND, VCC, GND_0, VCC_0;
    
    DFN1E1 \sd_sacq_data3[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[1]_net_1 ));
    NOR3A \i_RNO[6]  (.A(net_27), .B(N_577), .C(un1_i_reg18_1), .Y(
        \i_RNO[6]_net_1 ));
    XNOR2 \sd_sacq_data6_RNIGBB4[16]  (.A(count[16]), .B(
        \sd_sacq_data6[16]_net_1 ), .Y(N_371_i_i));
    DFN1E0 \sd_sacq_data5[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[2]_net_1 ));
    DFN1E0 \sd_sacq_data5[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[8]_net_1 ));
    NOR2B \i_RNO[2]  (.A(s_acq180_c), .B(net_27), .Y(\i_RNO_1[2] ));
    OR3C sd_sacq_data6_109_e (.A(N_573_1), .B(
        un1_sd_sacq_data117_1_i_a2_0), .C(sd_sacq_choice[0]), .Y(
        N_701_i));
    DFN1E1 \sd_sacq_data2[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[3]_net_1 ));
    DFN1 \i[7]  (.D(\i_RNO[7]_net_1 ), .CLK(ddsclkout_c), .Q(i[7]));
    DFN1E0 \sd_sacq_data4[20]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[20]_net_1 ));
    XNOR2 \sd_sacq_data1_RNI1G97[2]  (.A(count_4[2]), .B(
        \sd_sacq_data1[2]_net_1 ), .Y(N_420_i_i_0));
    DFN1E0 \sd_sacq_data6[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[7]_net_1 ));
    NOR3C \sd_sacq_data4_RNI8K7Q[15]  (.A(N_361_i_i), .B(N_337_i_i), 
        .C(\un1_count_NE_9[0] ), .Y(\un1_count_NE_15[0] ));
    DFN1E1 \sd_sacq_data2[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[4]_net_1 ));
    OR3A sd_sacq_data5_87_e (.A(sd_sacq_choice[0]), .B(N_580), .C(
        un1_sd_sacq_data117_2_i_a2_0_net_1), .Y(N_657));
    XA1A \sd_sacq_data1_RNI6MK8[13]  (.A(\sd_sacq_data1[13]_net_1 ), 
        .B(count[13]), .C(N_397_i_i_0), .Y(\i_reg18_NE_i_a2_2[0] ));
    DFN1E0 \sd_sacq_data6[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[12]_net_1 ));
    XNOR2 \sd_sacq_data4_RNI0G97[0]  (.A(count_4[0]), .B(
        \sd_sacq_data4[0]_net_1 ), .Y(N_357_i_i));
    DFN1E0 \sd_sacq_data4[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[11]_net_1 ));
    NOR2A un1_sd_sacq_data117_i_a2_0 (.A(sd_sacq_choice[1]), .B(
        sd_sacq_choice[2]), .Y(N_792));
    XA1A \sd_sacq_data2_RNIEEL8[12]  (.A(\sd_sacq_data2[12]_net_1 ), 
        .B(count[12]), .C(N_388_i_i_0), .Y(\un1_count_4_NE_i_a2_4[0] ));
    DFN1E1 \sd_sacq_data1[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[6]_net_1 ));
    DFN1E1 \sd_sacq_data1[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[1]_net_1 ));
    DFN1E1 \sd_sacq_data3[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[5]_net_1 ));
    DFN1E0 \sd_sacq_data7[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[0]_net_1 ));
    NOR3C \sd_sacq_data4_RNIIVHB2[3]  (.A(\un1_count_NE_11[0] ), .B(
        \un1_count_NE_10[0] ), .C(\un1_count_NE_17[0] ), .Y(
        \un1_count_NE_19[0] ));
    NOR3B sd_sacq_data1_0_sqmuxa_0_a2 (.A(sd_sacq_choice[0]), .B(
        un1_sd_sacq_data117_1_i_a2_0), .C(N_580), .Y(
        sd_sacq_data1_0_sqmuxa));
    DFN1E0 \sd_sacq_data5[20]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[20]_net_1 ));
    DFN1E0 \sd_sacq_data6[17]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[17]_net_1 ));
    NOR3C \sd_sacq_data4_RNIKPHB1[20]  (.A(\un1_count_NE_3[0] ), .B(
        \un1_count_NE_2[0] ), .C(\un1_count_NE_13[0] ), .Y(
        \un1_count_NE_17[0] ));
    DFN1 \i[0]  (.D(\i_RNO_1[0] ), .CLK(ddsclkout_c), .Q(i_4[0]));
    XNOR2 \sd_sacq_data4_RNIEG97[7]  (.A(count_1[7]), .B(
        \sd_sacq_data4[7]_net_1 ), .Y(N_305_i_i));
    NOR3C \sd_sacq_data3_RNI26GE1[12]  (.A(\un1_count_5_NE_i_a2_4[0] ), 
        .B(\un1_count_5_NE_i_a2_3[0] ), .C(\un1_count_5_NE_i_a2_9[0] ), 
        .Y(\un1_count_5_NE_i_a2_13[0] ));
    XA1A \sd_sacq_data1_RNIK0JE[8]  (.A(\sd_sacq_data1[8]_net_1 ), .B(
        count[8]), .C(N_378_i_i_0), .Y(\i_reg18_NE_i_a2_1[0] ));
    NOR2B \i_RNO[3]  (.A(scalestate_0_long_opentime), .B(net_27), .Y(
        \i_RNO_1[3] ));
    DFN1E0 \sd_sacq_data4[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[8]_net_1 ));
    DFN1E0 \sd_sacq_data5[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[4]_net_1 ));
    XNOR2 \i_RNO_17[10]  (.A(count[15]), .B(\sd_sacq_data7[15]_net_1 ), 
        .Y(N_340_i_i_0));
    XA1A \i_RNO_27[10]  (.A(\sd_sacq_data7[7]_net_1 ), .B(count_1[7]), 
        .C(N_324_i_i_0), .Y(\i_0_5[10] ));
    NOR3B \i_RNO[5]  (.A(net_27), .B(N_579), .C(N_578_i), .Y(
        \i_RNO[5]_net_1 ));
    XA1A \sd_sacq_data6_RNIU0JE[4]  (.A(\sd_sacq_data6[4]_net_1 ), .B(
        count_4[4]), .C(N_315_i_i), .Y(\un1_count_2_NE_9[0] ));
    NOR2A \i_RNO[4]  (.A(net_27), .B(N_579), .Y(\i_RNO[4]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIBRA4[14]  (.A(count[14]), .B(
        \sd_sacq_data5[14]_net_1 ), .Y(N_334_i_i));
    XNOR2 \sd_sacq_data2_RNI8G97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data2[5]_net_1 ), .Y(N_387_i_i_0));
    XA1A \sd_sacq_data6_RNI6FN8[19]  (.A(\sd_sacq_data6[19]_net_1 ), 
        .B(count[19]), .C(N_371_i_i), .Y(\un1_count_2_NE_1[0] ));
    XA1A \sd_sacq_data5_RNIOML8[21]  (.A(\sd_sacq_data5[21]_net_1 ), 
        .B(count[21]), .C(N_374_i_i), .Y(\un1_count_1_NE_0[0] ));
    XNOR2 \sd_sacq_data2_RNIAG97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data2[6]_net_1 ), .Y(N_395_i_i_0));
    OR2B \sd_sacq_data4_RNI7FHJF[10]  (.A(\un1_count_NE[0] ), .B(
        un1_count_6), .Y(un1_count_8));
    DFN1E0 \sd_sacq_data7[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[9]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIFBB4[16]  (.A(count[16]), .B(
        \sd_sacq_data5[16]_net_1 ), .Y(N_370_i_i));
    DFN1E1 \sd_sacq_data1[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[12]_net_1 ));
    DFN1E0 \sd_sacq_data4[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[1]_net_1 ));
    XNOR2 \sd_sacq_data4_RNIIRB4[18]  (.A(count[18]), .B(
        \sd_sacq_data4[18]_net_1 ), .Y(N_349_i_i));
    OR3A sd_sacq_data4_65_e (.A(sd_sacq_choice[0]), .B(N_580), .C(
        un1_sd_sacq_data117_3_i_a2_0_net_1), .Y(N_613));
    DFN1E0 \sd_sacq_data4[21]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[21]_net_1 ));
    XNOR2 \i_RNO_32[10]  (.A(count_4[2]), .B(\sd_sacq_data7[2]_net_1 ), 
        .Y(N_344_i_i_0));
    DFN1E0 \sd_sacq_data6[19]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[19]_net_1 ));
    XA1A \sd_sacq_data4_RNIQ0JE[4]  (.A(\sd_sacq_data4[4]_net_1 ), .B(
        count_4[4]), .C(N_313_i_i), .Y(\un1_count_NE_9[0] ));
    DFN1E0 \sd_sacq_data7[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[6]_net_1 ));
    XNOR2 \sd_sacq_data2_RNI23A4[11]  (.A(count[11]), .B(
        \sd_sacq_data2[11]_net_1 ), .Y(N_392_i_i_0));
    NOR2B \i_RNO_4[10]  (.A(N_360_i_i_0), .B(\i_0_0[10] ), .Y(
        \i_0_11[10] ));
    XA1A \sd_sacq_data6_RNIC6K8[10]  (.A(\sd_sacq_data6[10]_net_1 ), 
        .B(count[10]), .C(N_327_i_i), .Y(\un1_count_2_NE_7[0] ));
    XNOR2 \sd_sacq_data5_RNI3G97[1]  (.A(count_4[1]), .B(
        \sd_sacq_data5[1]_net_1 ), .Y(N_362_i_i));
    XNOR2 \sd_sacq_data4_RNIIG97[9]  (.A(count[9]), .B(
        \sd_sacq_data4[9]_net_1 ), .Y(N_313_i_i));
    DFN1E0 \sd_sacq_data6[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[15]_net_1 ));
    XA1A \sd_sacq_data2_RNI6BJB[10]  (.A(\sd_sacq_data2[10]_net_1 ), 
        .B(count[10]), .C(N_416_i_i_0), .Y(\un1_count_4_NE_i_a2_6[0] ));
    NOR3C \sd_sacq_data6_RNI4QHB1[18]  (.A(\un1_count_2_NE_3[0] ), .B(
        \un1_count_2_NE_2[0] ), .C(\un1_count_2_NE_13[0] ), .Y(
        \un1_count_2_NE_17[0] ));
    XNOR2 \sd_sacq_data4_RNI6BA4[12]  (.A(count[12]), .B(
        \sd_sacq_data4[12]_net_1 ), .Y(N_325_i_i));
    XNOR2 \sd_sacq_data4_RNIARA4[14]  (.A(count[14]), .B(
        \sd_sacq_data4[14]_net_1 ), .Y(N_333_i_i));
    XNOR2 \sd_sacq_data6_RNIIJB4[17]  (.A(count[17]), .B(
        \sd_sacq_data6[17]_net_1 ), .Y(N_375_i_i));
    DFN1E0 \sd_sacq_data6[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[13]_net_1 ));
    XNOR2 \sd_sacq_data3_RNI5G97[3]  (.A(count_4[3]), .B(
        \sd_sacq_data3[3]_net_1 ), .Y(N_384_i_i_0));
    XNOR2 \sd_sacq_data1_RNI9G97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data1[6]_net_1 ), .Y(N_400_i_i_0));
    DFN1E0 \sd_sacq_data5[21]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[21]_net_1 ));
    XNOR2 \i_RNO_31[10]  (.A(count[11]), .B(\sd_sacq_data7[11]_net_1 ), 
        .Y(N_324_i_i_0));
    DFN1E1 \sd_sacq_data2[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[9]_net_1 ));
    OR2B \sd_sacq_data2_RNIUNLP7[10]  (.A(N_579), .B(N_578_i), .Y(
        un1_i_reg18_1));
    XNOR2 \sd_sacq_data4_RNI8JA4[13]  (.A(count[13]), .B(
        \sd_sacq_data4[13]_net_1 ), .Y(N_329_i_i));
    NOR2B \i_RNO[0]  (.A(scalestate_0_s_acq), .B(net_27), .Y(
        \i_RNO_1[0] ));
    XA1A \sd_sacq_data5_RNISBKB[8]  (.A(\sd_sacq_data5[8]_net_1 ), .B(
        count[8]), .C(N_334_i_i), .Y(\un1_count_1_NE_2[0] ));
    XA1A \sd_sacq_data5_RNIOML8[18]  (.A(\sd_sacq_data5[18]_net_1 ), 
        .B(count[18]), .C(\un1_count_1_20_i[0] ), .Y(
        \un1_count_1_NE_3[0] ));
    NOR3C \sd_sacq_data5_RNI8N7N[11]  (.A(N_306_i_i), .B(N_294_i_i), 
        .C(\un1_count_1_NE_5[0] ), .Y(\un1_count_1_NE_13[0] ));
    XNOR2 \sd_sacq_data6_RNIE3B4[15]  (.A(count[15]), .B(
        \sd_sacq_data6[15]_net_1 ), .Y(N_339_i_i));
    OR2A un1_sd_sacq_data117_2_i_a2_0 (.A(top_code_0_sd_sacq_load), .B(
        sd_sacq_choice[3]), .Y(N_580));
    XNOR2 \sd_sacq_data6_RNI8BA4[12]  (.A(count[12]), .B(
        \sd_sacq_data6[12]_net_1 ), .Y(N_327_i_i));
    DFN1E0 \sd_sacq_data6[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[1]_net_1 ));
    NOR3C \sd_sacq_data2_RNI6SGU[0]  (.A(N_394_i_i_0), .B(N_389_i_i_0), 
        .C(\un1_count_4_NE_i_a2_8[0] ), .Y(\un1_count_4_NE_i_a2_12[0] )
        );
    XA1C \sd_sacq_data1_RNIJBK8[14]  (.A(\sd_sacq_data1[14]_net_1 ), 
        .B(count[14]), .C(count[20]), .Y(\i_reg18_NE_i_a2_0[0] ));
    GND GND_i (.Y(GND));
    DFN1E0 \sd_sacq_data6[18]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[18]_net_1 ));
    NOR2B \sd_sacq_data4_RNICMK8[11]  (.A(N_321_i_i), .B(N_329_i_i), 
        .Y(\un1_count_NE_5[0] ));
    XA1A \sd_sacq_data5_RNII0JE[2]  (.A(\sd_sacq_data5[2]_net_1 ), .B(
        count_4[2]), .C(N_302_i_i), .Y(\un1_count_1_NE_6[0] ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1E0 \sd_sacq_data7[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[4]_net_1 ));
    XA1A \sd_sacq_data2_RNIIRTF[0]  (.A(\sd_sacq_data2[0]_net_1 ), .B(
        count_4[0]), .C(\un1_count_4_NE_i_a2_0[0] ), .Y(
        \un1_count_4_NE_i_a2_8[0] ));
    XNOR2 \sd_sacq_data6_RNIAJA4[13]  (.A(count[13]), .B(
        \sd_sacq_data6[13]_net_1 ), .Y(N_331_i_i));
    NOR3C \i_RNO_8[10]  (.A(N_368_i_i_0), .B(N_364_i_i_0), .C(
        \i_0_10[10] ), .Y(\i_0_16[10] ));
    DFN1E1 \sd_sacq_data1[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[15]_net_1 ));
    DFN1E0 \sd_sacq_data6[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[10]_net_1 ));
    DFN1E1 \sd_sacq_data2[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[12]_net_1 ));
    DFN1E1 \sd_sacq_data1[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[13]_net_1 ));
    NOR2B \sd_sacq_data4_RNI2FN8[16]  (.A(N_353_i_i), .B(N_369_i_i), 
        .Y(\un1_count_NE_1[0] ));
    DFN1E0 \sd_sacq_data5[16]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[16]_net_1 ));
    XNOR2 \sd_sacq_data4_RNIK3C4[19]  (.A(count[19]), .B(
        \sd_sacq_data4[19]_net_1 ), .Y(N_353_i_i));
    XA1A \sd_sacq_data4_RNI60JE[3]  (.A(\sd_sacq_data4[3]_net_1 ), .B(
        count_4[3]), .C(N_357_i_i), .Y(\un1_count_NE_10[0] ));
    OR3C \sd_sacq_data1_RNINRQS3[10]  (.A(\i_reg18_NE_i_a2_13[0] ), .B(
        \i_reg18_NE_i_a2_12[0] ), .C(\i_reg18_NE_i_a2_14[0] ), .Y(
        N_579));
    NOR3C \i_RNO_1[10]  (.A(\i_0_12[10] ), .B(\i_0_11[10] ), .C(
        \i_0_18[10] ), .Y(\i_0_20[10] ));
    XNOR2 \sd_sacq_data4_RNIGJB4[17]  (.A(count[17]), .B(
        \sd_sacq_data4[17]_net_1 ), .Y(N_373_i_i));
    DFN1E0 \sd_sacq_data6[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[2]_net_1 ));
    OR3C sd_sacq_data7_131_e (.A(N_573_1), .B(N_792), .C(
        sd_sacq_choice[0]), .Y(N_745_i));
    XNOR2 \sd_sacq_data6_RNIEG97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data6[6]_net_1 ), .Y(N_303_i_i));
    DFN1E0 \sd_sacq_data5[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[7]_net_1 ));
    NOR2B \i_RNO_15[10]  (.A(\i_0_5[10] ), .B(\i_0_6[10] ), .Y(
        \i_0_14[10] ));
    NOR3C \sd_sacq_data5_RNI46001[21]  (.A(\un1_count_1_NE_1[0] ), .B(
        \un1_count_1_NE_0[0] ), .C(\un1_count_1_NE_10[0] ), .Y(
        \un1_count_1_NE_16[0] ));
    NOR2B un1_sd_sacq_data117_i_a2_1 (.A(sd_sacq_choice[3]), .B(
        top_code_0_sd_sacq_load), .Y(N_573_1));
    XNOR2 \i_RNO_25[10]  (.A(count_1[5]), .B(\sd_sacq_data7[5]_net_1 ), 
        .Y(N_296_i_i_0));
    DFN1 \i[9]  (.D(\i_RNO[9]_net_1 ), .CLK(ddsclkout_c), .Q(i[9]));
    XNOR2 \sd_sacq_data4_RNI63A4[21]  (.A(count[21]), .B(
        \sd_sacq_data4[21]_net_1 ), .Y(N_297_i_i));
    XA1A \sd_sacq_data6_RNIQML8[21]  (.A(\sd_sacq_data6[21]_net_1 ), 
        .B(count[21]), .C(N_375_i_i), .Y(\un1_count_2_NE_0[0] ));
    DFN1E0 \sd_sacq_data6[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[3]_net_1 ));
    DFN1E0 \sd_sacq_data5[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[5]_net_1 ));
    DFN1E0 \sd_sacq_data6[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[14]_net_1 ));
    DFN1E0 \sd_sacq_data4[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[6]_net_1 ));
    DFN1E1 \sd_sacq_data3[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[2]_net_1 ));
    XA1A \sd_sacq_data5_RNIS0JE[4]  (.A(\sd_sacq_data5[4]_net_1 ), .B(
        count_4[4]), .C(N_314_i_i), .Y(\un1_count_1_NE_9[0] ));
    NOR3A sd_sacq_data2_1_sqmuxa_0_a2 (.A(N_792), .B(sd_sacq_choice[0])
        , .C(N_580), .Y(sd_sacq_data2_1_sqmuxa));
    XNOR2 \sd_sacq_data4_RNI2G97[1]  (.A(count_4[1]), .B(
        \sd_sacq_data4[1]_net_1 ), .Y(N_361_i_i));
    DFN1E1 \sd_sacq_data3[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[6]_net_1 ));
    OR3C \sd_sacq_data2_RNI7SQS3[10]  (.A(\un1_count_4_NE_i_a2_13[0] ), 
        .B(\un1_count_4_NE_i_a2_12[0] ), .C(
        \un1_count_4_NE_i_a2_14[0] ), .Y(N_578_i));
    XNOR2 \sd_sacq_data2_RNICG97[7]  (.A(count_1[7]), .B(
        \sd_sacq_data2[7]_net_1 ), .Y(N_393_i_i_0));
    VCC VCC_i (.Y(VCC));
    DFN1E0 \sd_sacq_data5[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[12]_net_1 ));
    XNOR2 \sd_sacq_data3_RNIBG97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data3[6]_net_1 ), .Y(N_405_i_i_0));
    XA1A \i_RNO_9[10]  (.A(\sd_sacq_data7[17]_net_1 ), .B(count[17]), 
        .C(N_356_i_i_0), .Y(\i_0_1[10] ));
    XA1A \i_RNO_10[10]  (.A(\sd_sacq_data7[16]_net_1 ), .B(count[16]), 
        .C(N_312_i_i_0), .Y(\i_0_2[10] ));
    OR3 sd_sacq_data5_71_e (.A(N_580), .B(
        un1_sd_sacq_data117_2_i_a2_0_net_1), .C(sd_sacq_choice[0]), .Y(
        N_625_i));
    DFN1E0 \sd_sacq_data5[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[6]_net_1 ));
    DFN1E1 \sd_sacq_data2[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[7]_net_1 ));
    XNOR2 \i_RNO_20[10]  (.A(count_4[4]), .B(\sd_sacq_data7[4]_net_1 ), 
        .Y(N_368_i_i_0));
    XNOR2 \sd_sacq_data5_RNID3B4[15]  (.A(count[15]), .B(
        \sd_sacq_data5[15]_net_1 ), .Y(N_338_i_i));
    NOR2B \sd_sacq_data4_RNIQBKB[14]  (.A(N_309_i_i), .B(N_333_i_i), 
        .Y(\un1_count_NE_2[0] ));
    NOR3C \sd_sacq_data6_RNIGREH1[10]  (.A(\un1_count_2_NE_7[0] ), .B(
        \un1_count_2_NE_6[0] ), .C(\un1_count_2_NE_15[0] ), .Y(
        \un1_count_2_NE_18[0] ));
    DFN1E0 \sd_sacq_data6[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[5]_net_1 ));
    DFN1E1 \sd_sacq_data1[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[10]_net_1 ));
    OR2A \i_RNO_0[9]  (.A(net_27), .B(\un1_count_2_i[0] ), .Y(
        \i_0_0[9] ));
    DFN1E0 \sd_sacq_data5[17]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[17]_net_1 ));
    XA1A \sd_sacq_data3_RNIAMK8[13]  (.A(\sd_sacq_data3[13]_net_1 ), 
        .B(count[13]), .C(N_402_i_i_0), .Y(\un1_count_5_NE_i_a2_2[0] ));
    XNOR2 \sd_sacq_data5_RNIHJB4[17]  (.A(count[17]), .B(
        \sd_sacq_data5[17]_net_1 ), .Y(N_374_i_i));
    DFN1E1 \sd_sacq_data3[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[9]_net_1 ));
    DFN1E1 \sd_sacq_data3[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[4]_net_1 ));
    XNOR2 \sd_sacq_data2_RNI6G97[4]  (.A(count_4[4]), .B(
        \sd_sacq_data2[4]_net_1 ), .Y(N_416_i_i_0));
    OR3B sd_sacq_data6_100_e (.A(N_573_1), .B(
        un1_sd_sacq_data117_1_i_a2_0), .C(sd_sacq_choice[0]), .Y(
        N_683_i));
    DFN1E0 \sd_sacq_data4[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[0]_net_1 ));
    XNOR2 \sd_sacq_data3_RNI33A4[11]  (.A(count[11]), .B(
        \sd_sacq_data3[11]_net_1 ), .Y(N_402_i_i_0));
    XNOR2 \i_RNO_19[10]  (.A(count[10]), .B(\sd_sacq_data7[10]_net_1 ), 
        .Y(N_320_i_i_0));
    DFN1E0 \sd_sacq_data6[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[11]_net_1 ));
    XA1A \sd_sacq_data5_RNI80JE[3]  (.A(\sd_sacq_data5[3]_net_1 ), .B(
        count_4[3]), .C(N_358_i_i), .Y(\un1_count_1_NE_10[0] ));
    DFN1E1 \sd_sacq_data2[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[15]_net_1 ));
    XNOR2 \i_RNO_29[10]  (.A(count[9]), .B(\sd_sacq_data7[9]_net_1 ), 
        .Y(N_316_i_i_0));
    XA1A \sd_sacq_data3_RNIKRTF[0]  (.A(\sd_sacq_data3[0]_net_1 ), .B(
        count_4[0]), .C(\un1_count_5_NE_i_a2_0[0]_net_1 ), .Y(
        \un1_count_5_NE_i_a2_8[0] ));
    XA1A \sd_sacq_data5_RNIA6K8[10]  (.A(\sd_sacq_data5[10]_net_1 ), 
        .B(count[10]), .C(N_326_i_i), .Y(\un1_count_1_NE_7[0] ));
    DFN1E1 \sd_sacq_data2[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[13]_net_1 ));
    XA1A \sd_sacq_data6_RNIQML8[18]  (.A(\sd_sacq_data6[18]_net_1 ), 
        .B(count[18]), .C(\un1_count_2_20_i[0] ), .Y(
        \un1_count_2_NE_3[0] ));
    XNOR2 \sd_sacq_data2_RNIGG97[9]  (.A(count[9]), .B(
        \sd_sacq_data2[9]_net_1 ), .Y(N_394_i_i_0));
    DFN1E1 \sd_sacq_data3[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[12]_net_1 ));
    DFN1E1 \sd_sacq_data1[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[14]_net_1 ));
    XA1A \i_RNO_14[10]  (.A(\sd_sacq_data7[14]_net_1 ), .B(count[14]), 
        .C(N_352_i_i_0), .Y(\i_0_3[10] ));
    DFN1E0 \sd_sacq_data7[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[8]_net_1 ));
    NOR3C \sd_sacq_data4_RNI0REH1[10]  (.A(\un1_count_NE_7[0] ), .B(
        \un1_count_NE_6[0] ), .C(\un1_count_NE_15[0] ), .Y(
        \un1_count_NE_18[0] ));
    XNOR2 \i_RNO_24[10]  (.A(count[8]), .B(\sd_sacq_data7[8]_net_1 ), 
        .Y(N_312_i_i_0));
    NOR3A \i_RNO[9]  (.A(\un1_count_1_NE[0] ), .B(un1_count_8), .C(
        \i_0_0[9] ), .Y(\i_RNO[9]_net_1 ));
    DFN1E1 \sd_sacq_data2[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[2]_net_1 ));
    DFN1E1 \sd_sacq_data1[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[9]_net_1 ));
    NOR3C \sd_sacq_data6_RNICN7N[11]  (.A(N_307_i_i), .B(N_295_i_i), 
        .C(\un1_count_2_NE_5[0] ), .Y(\un1_count_2_NE_13[0] ));
    DFN1E0 \sd_sacq_data7[16]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[16]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIBG97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data5[5]_net_1 ), .Y(N_294_i_i));
    XNOR2 \sd_sacq_data4_RNIC3B4[15]  (.A(count[15]), .B(
        \sd_sacq_data4[15]_net_1 ), .Y(N_337_i_i));
    XNOR2 \sd_sacq_data1_RNI13A4[11]  (.A(count[11]), .B(
        \sd_sacq_data1[11]_net_1 ), .Y(N_397_i_i_0));
    DFN1E0 \sd_sacq_data5[19]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[19]_net_1 ));
    NOR3C \i_RNO_0[10]  (.A(\i_0_20[10] ), .B(\i_0_19[10] ), .C(
        \un1_count_2_i[0] ), .Y(\i_0_22[10] ));
    DFN1E0 \sd_sacq_data6[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[9]_net_1 ));
    XNOR2 \sd_sacq_data3_RNI9G97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data3[5]_net_1 ), .Y(N_383_i_i_0));
    DFN1E0 \sd_sacq_data5[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[15]_net_1 ));
    NOR3C \sd_sacq_data3_RNI2N7N[13]  (.A(N_383_i_i_0), .B(N_409_i_i_0)
        , .C(\un1_count_5_NE_i_a2_2[0] ), .Y(
        \un1_count_5_NE_i_a2_9[0] ));
    DFN1E1 \sd_sacq_data1[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[7]_net_1 ));
    NOR3C \sd_sacq_data3_RNIASGU[0]  (.A(N_404_i_i_0), .B(N_384_i_i_0), 
        .C(\un1_count_5_NE_i_a2_8[0] ), .Y(\un1_count_5_NE_i_a2_12[0] )
        );
    XNOR2 \sd_sacq_data1_RNIFG97[9]  (.A(count[9]), .B(
        \sd_sacq_data1[9]_net_1 ), .Y(N_399_i_i_0));
    DFN1E1 \sd_sacq_data1[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[3]_net_1 ));
    DFN1E0 \sd_sacq_data5[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[13]_net_1 ));
    NOR3B sd_sacq_data3_1_sqmuxa_0_a2 (.A(N_792), .B(sd_sacq_choice[0])
        , .C(N_580), .Y(sd_sacq_data3_1_sqmuxa));
    DFN1E1 \sd_sacq_data1[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[11]_net_1 ));
    OR2B un1_sd_sacq_data117_2_i_a2_0_0 (.A(sd_sacq_choice[1]), .B(
        sd_sacq_choice[2]), .Y(un1_sd_sacq_data117_2_i_a2_0_net_1));
    XNOR2 \sd_sacq_data4_RNIGG97[8]  (.A(count[8]), .B(
        \sd_sacq_data4[8]_net_1 ), .Y(N_309_i_i));
    DFN1 \i[2]  (.D(\i_RNO_1[2] ), .CLK(ddsclkout_c), .Q(i_3[2]));
    DFN1E1 \sd_sacq_data2[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[10]_net_1 ));
    DFN1E0 \sd_sacq_data7[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[12]_net_1 ));
    OR3 sd_sacq_data4_49_e (.A(N_580), .B(
        un1_sd_sacq_data117_3_i_a2_0_net_1), .C(sd_sacq_choice[0]), .Y(
        N_581_i));
    DFN1E1 \sd_sacq_data1[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[0]_net_1 ));
    XNOR2 \sd_sacq_data5_RNI1G97[0]  (.A(count_4[0]), .B(
        \sd_sacq_data5[0]_net_1 ), .Y(N_358_i_i));
    DFN1E1 \sd_sacq_data1[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[5]_net_1 ));
    XA1A \i_RNO_13[10]  (.A(\sd_sacq_data7[20]_net_1 ), .B(count[20]), 
        .C(N_296_i_i_0), .Y(\i_0_4[10] ));
    XNOR2 \i_RNO_23[10]  (.A(count[19]), .B(\sd_sacq_data7[19]_net_1 ), 
        .Y(N_356_i_i_0));
    DFN1E1 \sd_sacq_data2[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[8]_net_1 ));
    DFN1E0 \sd_sacq_data7[17]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[17]_net_1 ));
    XA1A \sd_sacq_data6_RNIK0JE[2]  (.A(\sd_sacq_data6[2]_net_1 ), .B(
        count_4[2]), .C(N_303_i_i), .Y(\un1_count_2_NE_6[0] ));
    XA1A \sd_sacq_data1_RNIGRTF[0]  (.A(\sd_sacq_data1[0]_net_1 ), .B(
        count_4[0]), .C(\i_reg18_NE_i_a2_0[0] ), .Y(
        \i_reg18_NE_i_a2_8[0] ));
    DFN1E0 \sd_sacq_data5[18]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_657), .Q(\sd_sacq_data5[18]_net_1 ));
    XNOR2 \sd_sacq_data4_RNIEBB4[16]  (.A(count[16]), .B(
        \sd_sacq_data4[16]_net_1 ), .Y(N_369_i_i));
    DFN1E0 \sd_sacq_data7[20]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[20]_net_1 ));
    DFN1E1 \sd_sacq_data3[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[15]_net_1 ));
    NOR3C \sd_sacq_data1_RNI3QPF1[10]  (.A(\i_reg18_NE_i_a2_6[0] ), .B(
        \i_reg18_NE_i_a2_5[0] ), .C(N_904), .Y(\i_reg18_NE_i_a2_14[0] )
        );
    XA1A \i_RNO_12[10]  (.A(\sd_sacq_data7[21]_net_1 ), .B(count[21]), 
        .C(net_27), .Y(\i_0_0[10] ));
    NOR2B \i_RNO_3[10]  (.A(\i_0_1[10] ), .B(\i_0_2[10] ), .Y(
        \i_0_12[10] ));
    NOR2B \i_RNO_22[10]  (.A(N_316_i_i_0), .B(N_348_i_i_0), .Y(
        \i_0_10[10] ));
    NOR3A \un1_count_5_NE_i_a2_0[0]  (.A(
        \un1_count_5_NE_i_a2_0_2[0]_net_1 ), .B(count[19]), .C(
        count[16]), .Y(N_904));
    DFN1E1 \sd_sacq_data3[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[13]_net_1 ));
    DFN1E1 \sd_sacq_data2[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[14]_net_1 ));
    DFN1 \i[10]  (.D(\i_RNO[10]_net_1 ), .CLK(ddsclkout_c), .Q(i[10]));
    DFN1E0 \sd_sacq_data4[16]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[16]_net_1 ));
    XA1A \sd_sacq_data5_RNIEMK8[11]  (.A(\sd_sacq_data5[11]_net_1 ), 
        .B(count[11]), .C(N_330_i_i), .Y(\un1_count_1_NE_5[0] ));
    XA1A \sd_sacq_data4_RNIG0JE[2]  (.A(\sd_sacq_data4[2]_net_1 ), .B(
        count_4[2]), .C(N_301_i_i), .Y(\un1_count_NE_6[0] ));
    DFN1 \i[6]  (.D(\i_RNO[6]_net_1 ), .CLK(ddsclkout_c), .Q(i[6]));
    DFN1E1 \sd_sacq_data3[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[0]_net_1 ));
    DFN1E0 \sd_sacq_data4[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[4]_net_1 ));
    XNOR2 \sd_sacq_data5_RNI5R94[20]  (.A(count[20]), .B(
        \sd_sacq_data5[20]_net_1 ), .Y(\un1_count_1_20_i[0] ));
    DFN1 \i[4]  (.D(\i_RNO[4]_net_1 ), .CLK(ddsclkout_c), .Q(i[4]));
    DFN1E0 \sd_sacq_data5[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[10]_net_1 ));
    NOR2A \sd_sacq_data3_RNILKGMB[10]  (.A(N_577), .B(un1_i_reg18_1), 
        .Y(un1_count_6));
    XNOR2 \i_RNO_11[10]  (.A(count_4[0]), .B(\sd_sacq_data7[0]_net_1 ), 
        .Y(N_360_i_i_0));
    XNOR2 \i_RNO_21[10]  (.A(count_4[1]), .B(\sd_sacq_data7[1]_net_1 ), 
        .Y(N_364_i_i_0));
    NOR2B \sd_sacq_data4_RNIMML8[20]  (.A(N_349_i_i), .B(
        \un1_count_20_i[0] ), .Y(\un1_count_NE_3[0] ));
    XA1A \sd_sacq_data3_RNI8BJB[10]  (.A(\sd_sacq_data3[10]_net_1 ), 
        .B(count[10]), .C(N_411_i_i_0), .Y(\un1_count_5_NE_i_a2_6[0] ));
    NOR3C \sd_sacq_data1_RNII5GE1[13]  (.A(\i_reg18_NE_i_a2_2[0] ), .B(
        \i_reg18_NE_i_a2_1[0] ), .C(\i_reg18_NE_i_a2_10[0] ), .Y(
        \i_reg18_NE_i_a2_13[0] ));
    DFN1E0 \sd_sacq_data7[19]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[19]_net_1 ));
    XNOR2 \sd_sacq_data4_RNI43A4[11]  (.A(count[11]), .B(
        \sd_sacq_data4[11]_net_1 ), .Y(N_321_i_i));
    XNOR2 \sd_sacq_data3_RNIB3B4[15]  (.A(count[15]), .B(
        \sd_sacq_data3[15]_net_1 ), .Y(N_382_i_i_0));
    GND GND_i_0 (.Y(GND_0));
    OR3C \sd_sacq_data6_RNIUR0T3[10]  (.A(\un1_count_2_NE_17[0] ), .B(
        \un1_count_2_NE_16[0] ), .C(\un1_count_2_NE_18[0] ), .Y(
        \un1_count_2_i[0] ));
    DFN1E0 \sd_sacq_data4[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[5]_net_1 ));
    XA1C \sd_sacq_data2_RNIKBK8[14]  (.A(\sd_sacq_data2[14]_net_1 ), 
        .B(count[14]), .C(count[20]), .Y(\un1_count_4_NE_i_a2_0[0] ));
    XNOR2 \sd_sacq_data2_RNI4G97[3]  (.A(count_4[3]), .B(
        \sd_sacq_data2[3]_net_1 ), .Y(N_389_i_i_0));
    XA1A \sd_sacq_data6_RNIA0JE[3]  (.A(\sd_sacq_data6[3]_net_1 ), .B(
        count_4[3]), .C(N_359_i_i), .Y(\un1_count_2_NE_10[0] ));
    DFN1E0 \sd_sacq_data4[12]  (.D(sd_sacq_data[12]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[12]_net_1 ));
    OR2A un1_sd_sacq_data117_3_i_a2_0 (.A(sd_sacq_choice[2]), .B(
        sd_sacq_choice[1]), .Y(un1_sd_sacq_data117_3_i_a2_0_net_1));
    DFN1E1 \sd_sacq_data2[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[11]_net_1 ));
    DFN1E0 \sd_sacq_data7[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[15]_net_1 ));
    DFN1E0 \sd_sacq_data6[20]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[20]_net_1 ));
    DFN1E0 \sd_sacq_data5[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[14]_net_1 ));
    XNOR2 \sd_sacq_data4_RNI4R94[20]  (.A(count[20]), .B(
        \sd_sacq_data4[20]_net_1 ), .Y(\un1_count_20_i[0] ));
    XNOR2 \sd_sacq_data6_RNICG97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data6[5]_net_1 ), .Y(N_295_i_i));
    NOR3C \sd_sacq_data5_RNISPHB1[18]  (.A(\un1_count_1_NE_3[0] ), .B(
        \un1_count_1_NE_2[0] ), .C(\un1_count_1_NE_13[0] ), .Y(
        \un1_count_1_NE_17[0] ));
    XNOR2 \sd_sacq_data6_RNICRA4[14]  (.A(count[14]), .B(
        \sd_sacq_data6[14]_net_1 ), .Y(N_335_i_i));
    XNOR2 \sd_sacq_data4_RNICG97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data4[6]_net_1 ), .Y(N_301_i_i));
    XNOR2 \sd_sacq_data3_RNIHG97[9]  (.A(count[9]), .B(
        \sd_sacq_data3[9]_net_1 ), .Y(N_404_i_i_0));
    DFN1E0 \sd_sacq_data7[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[13]_net_1 ));
    NOR3C \sd_sacq_data5_RNI8REH1[10]  (.A(\un1_count_1_NE_7[0] ), .B(
        \un1_count_1_NE_6[0] ), .C(\un1_count_1_NE_15[0] ), .Y(
        \un1_count_1_NE_18[0] ));
    XNOR2 \i_RNO_18[10]  (.A(count_1[6]), .B(\sd_sacq_data7[6]_net_1 ), 
        .Y(N_304_i_i_0));
    OR3B sd_sacq_data7_115_e (.A(N_573_1), .B(N_792), .C(
        sd_sacq_choice[0]), .Y(N_713_i));
    DFN1E1 \sd_sacq_data3[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[10]_net_1 ));
    XNOR2 \sd_sacq_data6_RNI4G97[1]  (.A(count_4[1]), .B(
        \sd_sacq_data6[1]_net_1 ), .Y(N_363_i_i));
    DFN1E0 \sd_sacq_data4[17]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[17]_net_1 ));
    NOR3C \sd_sacq_data3_RNIBQPF1[10]  (.A(\un1_count_5_NE_i_a2_6[0] ), 
        .B(\un1_count_5_NE_i_a2_5[0] ), .C(N_904), .Y(
        \un1_count_5_NE_i_a2_14[0] ));
    XA1A \i_RNO_28[10]  (.A(\sd_sacq_data7[13]_net_1 ), .B(count[13]), 
        .C(N_344_i_i_0), .Y(\i_0_6[10] ));
    NOR3B \i_RNO[10]  (.A(\un1_count_1_NE[0] ), .B(\i_0_22[10] ), .C(
        un1_count_8), .Y(\i_RNO[10]_net_1 ));
    XNOR2 \sd_sacq_data2_RNIA3B4[15]  (.A(count[15]), .B(
        \sd_sacq_data2[15]_net_1 ), .Y(N_388_i_i_0));
    DFN1E1 \sd_sacq_data3[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[8]_net_1 ));
    DFN1E0 \sd_sacq_data7[21]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[21]_net_1 ));
    DFN1E1 \sd_sacq_data2[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[5]_net_1 ));
    NOR3C \i_RNO_5[10]  (.A(\i_0_4[10] ), .B(\i_0_3[10] ), .C(
        \i_0_14[10] ), .Y(\i_0_18[10] ));
    NOR3C \sd_sacq_data2_RNI7QPF1[10]  (.A(\un1_count_4_NE_i_a2_6[0] ), 
        .B(\un1_count_4_NE_i_a2_5[0] ), .C(N_904), .Y(
        \un1_count_4_NE_i_a2_14[0] ));
    DFN1E0 \sd_sacq_data5[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[3]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIDG97[6]  (.A(count_1[6]), .B(
        \sd_sacq_data5[6]_net_1 ), .Y(N_302_i_i));
    XA1A \sd_sacq_data5_RNI4FN8[19]  (.A(\sd_sacq_data5[19]_net_1 ), 
        .B(count[19]), .C(N_370_i_i), .Y(\un1_count_1_NE_1[0] ));
    XA1A \sd_sacq_data4_RNI86K8[10]  (.A(\sd_sacq_data4[10]_net_1 ), 
        .B(count[10]), .C(N_325_i_i), .Y(\un1_count_NE_7[0] ));
    XA1A \sd_sacq_data3_RNIC0JE[1]  (.A(\sd_sacq_data3[1]_net_1 ), .B(
        count_4[1]), .C(N_405_i_i_0), .Y(\un1_count_5_NE_i_a2_5[0] ));
    DFN1E1 \sd_sacq_data1[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[8]_net_1 ));
    NOR3A \i_RNO[8]  (.A(net_27), .B(\un1_count_1_NE[0] ), .C(
        un1_count_8), .Y(\i_RNO[8]_net_1 ));
    XNOR2 \sd_sacq_data1_RNI7G97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data1[5]_net_1 ), .Y(N_378_i_i_0));
    DFN1E0 \sd_sacq_data7[18]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_745_i), .Q(\sd_sacq_data7[18]_net_1 ));
    NOR3C \sd_sacq_data1_RNI2SGU[0]  (.A(N_399_i_i_0), .B(N_379_i_i_0), 
        .C(\i_reg18_NE_i_a2_8[0] ), .Y(\i_reg18_NE_i_a2_12[0] ));
    DFN1E1 \sd_sacq_data3[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[14]_net_1 ));
    DFN1E0 \sd_sacq_data4[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[2]_net_1 ));
    DFN1E0 \sd_sacq_data5[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[11]_net_1 ));
    DFN1E1 \sd_sacq_data3[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[3]_net_1 ));
    NOR3C \sd_sacq_data5_RNICK7Q[15]  (.A(N_362_i_i), .B(N_338_i_i), 
        .C(\un1_count_1_NE_9[0] ), .Y(\un1_count_1_NE_15[0] ));
    DFN1E1 \sd_sacq_data2[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[1]_net_1 ));
    XNOR2 \sd_sacq_data3_RNI3G97[2]  (.A(count_4[2]), .B(
        \sd_sacq_data3[2]_net_1 ), .Y(N_410_i_i_0));
    XA1A \sd_sacq_data6_RNIUBKB[8]  (.A(\sd_sacq_data6[8]_net_1 ), .B(
        count[8]), .C(N_335_i_i), .Y(\un1_count_2_NE_2[0] ));
    XA1A \sd_sacq_data2_RNIA0JE[1]  (.A(\sd_sacq_data2[1]_net_1 ), .B(
        count_4[1]), .C(N_395_i_i_0), .Y(\un1_count_4_NE_i_a2_5[0] ));
    NOR3C \sd_sacq_data1_RNIOE8N[12]  (.A(N_420_i_i_0), .B(N_398_i_i_0)
        , .C(\i_reg18_NE_i_a2_4[0] ), .Y(\i_reg18_NE_i_a2_10[0] ));
    NOR2 sd_sacq_data1_0_sqmuxa_0_a2_0 (.A(sd_sacq_choice[2]), .B(
        sd_sacq_choice[1]), .Y(un1_sd_sacq_data117_1_i_a2_0));
    XA1C \sd_sacq_data3_RNILBK8[14]  (.A(\sd_sacq_data3[14]_net_1 ), 
        .B(count[14]), .C(count[20]), .Y(
        \un1_count_5_NE_i_a2_0[0]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIJG97[9]  (.A(count[9]), .B(
        \sd_sacq_data5[9]_net_1 ), .Y(N_314_i_i));
    DFN1E0 \sd_sacq_data4[19]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[19]_net_1 ));
    XNOR2 \sd_sacq_data1_RNIBG97[7]  (.A(count_1[7]), .B(
        \sd_sacq_data1[7]_net_1 ), .Y(N_398_i_i_0));
    XNOR2 \sd_sacq_data1_RNI5G97[4]  (.A(count_4[4]), .B(
        \sd_sacq_data1[4]_net_1 ), .Y(N_421_i_i_0));
    DFN1E1 \sd_sacq_data1[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[2]_net_1 ));
    DFN1 \i[5]  (.D(\i_RNO[5]_net_1 ), .CLK(ddsclkout_c), .Q(i[5]));
    DFN1E0 \sd_sacq_data7[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[10]_net_1 ));
    XNOR2 \sd_sacq_data6_RNIGG97[7]  (.A(count_1[7]), .B(
        \sd_sacq_data6[7]_net_1 ), .Y(N_307_i_i));
    NOR3C \sd_sacq_data6_RNIA6001[21]  (.A(\un1_count_2_NE_1[0] ), .B(
        \un1_count_2_NE_0[0] ), .C(\un1_count_2_NE_10[0] ), .Y(
        \un1_count_2_NE_16[0] ));
    XA1A \sd_sacq_data2_RNI8MK8[13]  (.A(\sd_sacq_data2[13]_net_1 ), 
        .B(count[13]), .C(N_392_i_i_0), .Y(\un1_count_4_NE_i_a2_2[0] ));
    DFN1 \i[8]  (.D(\i_RNO[8]_net_1 ), .CLK(ddsclkout_c), .Q(i[8]));
    NOR3 \un1_count_5_NE_i_a2_0_2[0]  (.A(count[17]), .B(count[21]), 
        .C(count[18]), .Y(\un1_count_5_NE_i_a2_0_2[0]_net_1 ));
    XA1A \sd_sacq_data3_RNIG0JE[7]  (.A(\sd_sacq_data3[7]_net_1 ), .B(
        count_1[7]), .C(N_410_i_i_0), .Y(\un1_count_5_NE_i_a2_3[0] ));
    NOR2B \i_RNO_7[10]  (.A(N_304_i_i_0), .B(N_320_i_i_0), .Y(
        \i_0_7[10] ));
    DFN1E0 \sd_sacq_data4[15]  (.D(sd_sacq_data[15]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[15]_net_1 ));
    DFN1E0 \sd_sacq_data6[21]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[21]_net_1 ));
    XNOR2 \sd_sacq_data3_RNIFG97[8]  (.A(count[8]), .B(
        \sd_sacq_data3[8]_net_1 ), .Y(N_409_i_i_0));
    DFN1E0 \sd_sacq_data4[13]  (.D(sd_sacq_data[13]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[13]_net_1 ));
    NOR3C \sd_sacq_data4_RNIO5DH[21]  (.A(N_373_i_i), .B(N_297_i_i), 
        .C(\un1_count_NE_1[0] ), .Y(\un1_count_NE_11[0] ));
    DFN1E1 \sd_sacq_data3[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[11]_net_1 ));
    DFN1E0 \sd_sacq_data7[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[7]_net_1 ));
    XNOR2 \sd_sacq_data6_RNI2G97[0]  (.A(count_4[0]), .B(
        \sd_sacq_data6[0]_net_1 ), .Y(N_359_i_i));
    DFN1E0 \sd_sacq_data4[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[9]_net_1 ));
    DFN1E0 \sd_sacq_data7[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[14]_net_1 ));
    DFN1E1 \sd_sacq_data2[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[6]_net_1 ));
    NOR3C \i_RNO_2[10]  (.A(\i_0_8[10] ), .B(\i_0_7[10] ), .C(
        \i_0_16[10] ), .Y(\i_0_19[10] ));
    DFN1E0 \sd_sacq_data4[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[3]_net_1 ));
    DFN1E0 \sd_sacq_data4[18]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_613), .Q(\sd_sacq_data4[18]_net_1 ));
    DFN1 \i[3]  (.D(\i_RNO_1[3] ), .CLK(ddsclkout_c), .Q(i_3[3]));
    DFN1E1 \sd_sacq_data2[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        sd_sacq_data2_1_sqmuxa), .Q(\sd_sacq_data2[0]_net_1 ));
    NOR2B \i_RNO_6[10]  (.A(N_328_i_i_0), .B(N_340_i_i_0), .Y(
        \i_0_8[10] ));
    XA1A \sd_sacq_data6_RNIGMK8[11]  (.A(\sd_sacq_data6[11]_net_1 ), 
        .B(count[11]), .C(N_331_i_i), .Y(\un1_count_2_NE_5[0] ));
    OR3C \sd_sacq_data5_RNI8R0T3[10]  (.A(\un1_count_1_NE_17[0] ), .B(
        \un1_count_1_NE_16[0] ), .C(\un1_count_1_NE_18[0] ), .Y(
        \un1_count_1_NE[0] ));
    XA1A \sd_sacq_data2_RNIM0JE[8]  (.A(\sd_sacq_data2[8]_net_1 ), .B(
        count[8]), .C(N_387_i_i_0), .Y(\un1_count_4_NE_i_a2_1[0] ));
    DFN1E0 \sd_sacq_data7[3]  (.D(sd_sacq_data[3]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[3]_net_1 ));
    NOR3C \sd_sacq_data4_RNI4N7N[5]  (.A(N_305_i_i), .B(N_293_i_i), .C(
        \un1_count_NE_5[0] ), .Y(\un1_count_NE_13[0] ));
    NOR3C \sd_sacq_data2_RNIQ5GE1[13]  (.A(\un1_count_4_NE_i_a2_2[0] ), 
        .B(\un1_count_4_NE_i_a2_1[0] ), .C(\un1_count_4_NE_i_a2_10[0] )
        , .Y(\un1_count_4_NE_i_a2_13[0] ));
    DFN1E0 \sd_sacq_data6[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[4]_net_1 ));
    DFN1E0 \sd_sacq_data6[8]  (.D(sd_sacq_data[8]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[8]_net_1 ));
    NOR3C \sd_sacq_data6_RNIGK7Q[15]  (.A(N_363_i_i), .B(N_339_i_i), 
        .C(\un1_count_2_NE_9[0] ), .Y(\un1_count_2_NE_15[0] ));
    OR2B \sd_sacq_data4_RNIIQ0T3[10]  (.A(\un1_count_NE_19[0] ), .B(
        \un1_count_NE_18[0] ), .Y(\un1_count_NE[0] ));
    XNOR2 \sd_sacq_data6_RNI6R94[20]  (.A(count[20]), .B(
        \sd_sacq_data6[20]_net_1 ), .Y(\un1_count_2_20_i[0] ));
    DFN1E1 \sd_sacq_data3[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        sd_sacq_data3_1_sqmuxa), .Q(\sd_sacq_data3[7]_net_1 ));
    XA1A \sd_sacq_data1_RNI80JE[1]  (.A(\sd_sacq_data1[1]_net_1 ), .B(
        count_4[1]), .C(N_400_i_i_0), .Y(\i_reg18_NE_i_a2_5[0] ));
    XNOR2 \sd_sacq_data5_RNI7BA4[12]  (.A(count[12]), .B(
        \sd_sacq_data5[12]_net_1 ), .Y(N_326_i_i));
    DFN1 \i[1]  (.D(i_0_0_0), .CLK(ddsclkout_c), .Q(i_4[1]));
    DFN1E0 \sd_sacq_data7[2]  (.D(sd_sacq_data[2]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[2]_net_1 ));
    DFN1E0 \sd_sacq_data4[10]  (.D(sd_sacq_data[10]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[10]_net_1 ));
    NOR3B \i_RNO[7]  (.A(net_27), .B(un1_count_6), .C(
        \un1_count_NE[0] ), .Y(\i_RNO[7]_net_1 ));
    DFN1E0 \sd_sacq_data5[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[0]_net_1 ));
    DFN1E0 \sd_sacq_data7[11]  (.D(sd_sacq_data[11]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[11]_net_1 ));
    DFN1E0 \sd_sacq_data5[9]  (.D(sd_sacq_data[9]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[9]_net_1 ));
    XA1A \sd_sacq_data1_RNICEL8[12]  (.A(\sd_sacq_data1[12]_net_1 ), 
        .B(count[12]), .C(N_377_i_i_0), .Y(\i_reg18_NE_i_a2_4[0] ));
    XA1A \sd_sacq_data1_RNI4BJB[10]  (.A(\sd_sacq_data1[10]_net_1 ), 
        .B(count[10]), .C(N_421_i_i_0), .Y(\i_reg18_NE_i_a2_6[0] ));
    DFN1E0 \sd_sacq_data6[6]  (.D(sd_sacq_data[6]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[6]_net_1 ));
    XNOR2 \sd_sacq_data4_RNIAG97[5]  (.A(count_1[5]), .B(
        \sd_sacq_data4[5]_net_1 ), .Y(N_293_i_i));
    XNOR2 \sd_sacq_data5_RNI9JA4[13]  (.A(count[13]), .B(
        \sd_sacq_data5[13]_net_1 ), .Y(N_330_i_i));
    XA1A \sd_sacq_data3_RNIGEL8[12]  (.A(\sd_sacq_data3[12]_net_1 ), 
        .B(count[12]), .C(N_382_i_i_0), .Y(\un1_count_5_NE_i_a2_4[0] ));
    XNOR2 \i_RNO_30[10]  (.A(count_4[3]), .B(\sd_sacq_data7[3]_net_1 ), 
        .Y(N_348_i_i_0));
    NOR3C \sd_sacq_data2_RNISE8N[12]  (.A(N_415_i_i_0), .B(N_393_i_i_0)
        , .C(\un1_count_4_NE_i_a2_4[0] ), .Y(
        \un1_count_4_NE_i_a2_10[0] ));
    DFN1E1 \sd_sacq_data1[4]  (.D(sd_sacq_data[4]), .CLK(GLA), .E(
        sd_sacq_data1_0_sqmuxa), .Q(\sd_sacq_data1[4]_net_1 ));
    XNOR2 \sd_sacq_data3_RNI7G97[4]  (.A(count_4[4]), .B(
        \sd_sacq_data3[4]_net_1 ), .Y(N_411_i_i_0));
    DFN1E0 \sd_sacq_data5[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_625_i), .Q(\sd_sacq_data5[1]_net_1 ));
    XNOR2 \sd_sacq_data1_RNI3G97[3]  (.A(count_4[3]), .B(
        \sd_sacq_data1[3]_net_1 ), .Y(N_379_i_i_0));
    DFN1E0 \sd_sacq_data6[0]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_683_i), .Q(\sd_sacq_data6[0]_net_1 ));
    OR3C \sd_sacq_data3_RNINSQS3[10]  (.A(\un1_count_5_NE_i_a2_13[0] ), 
        .B(\un1_count_5_NE_i_a2_12[0] ), .C(
        \un1_count_5_NE_i_a2_14[0] ), .Y(N_577));
    DFN1E0 \sd_sacq_data7[1]  (.D(sd_sacq_data[1]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[1]_net_1 ));
    DFN1E0 \sd_sacq_data4[14]  (.D(sd_sacq_data[14]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[14]_net_1 ));
    DFN1E0 \sd_sacq_data6[16]  (.D(sd_sacq_data[0]), .CLK(GLA), .E(
        N_701_i), .Q(\sd_sacq_data6[16]_net_1 ));
    XNOR2 \i_RNO_16[10]  (.A(count[12]), .B(\sd_sacq_data7[12]_net_1 ), 
        .Y(N_328_i_i_0));
    DFN1E0 \sd_sacq_data7[5]  (.D(sd_sacq_data[5]), .CLK(GLA), .E(
        N_713_i), .Q(\sd_sacq_data7[5]_net_1 ));
    XNOR2 \sd_sacq_data5_RNIFG97[7]  (.A(count_1[7]), .B(
        \sd_sacq_data5[7]_net_1 ), .Y(N_306_i_i));
    XNOR2 \sd_sacq_data2_RNI2G97[2]  (.A(count_4[2]), .B(
        \sd_sacq_data2[2]_net_1 ), .Y(N_415_i_i_0));
    XNOR2 \sd_sacq_data1_RNI93B4[15]  (.A(count[15]), .B(
        \sd_sacq_data1[15]_net_1 ), .Y(N_377_i_i_0));
    XNOR2 \i_RNO_26[10]  (.A(count[18]), .B(\sd_sacq_data7[18]_net_1 ), 
        .Y(N_352_i_i_0));
    DFN1E0 \sd_sacq_data4[7]  (.D(sd_sacq_data[7]), .CLK(GLA), .E(
        N_581_i), .Q(\sd_sacq_data4[7]_net_1 ));
    XNOR2 \sd_sacq_data6_RNIKG97[9]  (.A(count[9]), .B(
        \sd_sacq_data6[9]_net_1 ), .Y(N_315_i_i));
    
endmodule


module sd_sacq_state(
       i_3,
       i_4,
       i,
       ddsclkout_c,
       sd_acq_en_c,
       sd_sacq_state_0_stateover,
       net_27
    );
input  [3:2] i_3;
input  [1:0] i_4;
input  [10:4] i;
input  ddsclkout_c;
output sd_acq_en_c;
output sd_sacq_state_0_stateover;
input  net_27;

    wire \cs_srsts_0_i_0[9] , \cs[5]_net_1 , cs4, \cs_srsts_0_i_0[12] , 
        en2_0_0_o3_0, N_201, N_232, N_233, ns_0_1_i_a2_1, 
        \cs[14]_net_1 , \cs[15]_net_1 , ns_0_1_i_a2_0, \cs[4]_net_1 , 
        \cs[11]_net_1 , N_245, \cs_RNO[14]_net_1 , \cs[13]_net_1 , 
        N_187_i_0, \cs_RNO_0[12]_net_1 , \cs[12]_net_1 , 
        \cs_RNO_0[11] , \cs[10]_net_1 , N_182_i_0, N_207, 
        \cs[9]_net_1 , \cs_RNO_1[6]_net_1 , N_218, N_219, 
        \cs_RNO_0[2]_net_1 , N_214, N_215, \cs_RNO_1[4] , en1, 
        \cs_RNO_2[5] , N_216, N_217, \cs_RNO_0[8]_net_1 , N_221, N_222, 
        \cs_RNO_2[3] , N_237, N_236, \cs[6]_net_1 , \cs_nsss[7] , 
        N_203, \cs_nsss[10] , \cs_nsss[13] , en2_RNO_net_1, N_230, 
        N_231, \cs_RNO_1[1] , \cs_i[0]_net_1 , \cs_RNO[15]_net_1 , 
        stateover_RNO_0, N_235, N_234, \cs[2]_net_1 , \cs[7]_net_1 , 
        \cs[8]_net_1 , \cs[1]_net_1 , en2_net_1, GND, VCC, GND_0, 
        VCC_0;
    
    NOR2 \cs_RNIT97E[6]  (.A(N_235), .B(N_234), .Y(N_203));
    NOR2A \cs_RNO[13]  (.A(cs4), .B(N_201), .Y(\cs_nsss[13] ));
    OA1 \cs_RNO[10]  (.A(N_232), .B(N_233), .C(cs4), .Y(\cs_nsss[10] ));
    DFN1 \cs[6]  (.D(\cs_RNO_1[6]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[6]_net_1 ));
    NOR2B \cs_RNI3V37[9]  (.A(i[7]), .B(\cs[9]_net_1 ), .Y(N_232));
    NOR3C \cs_RNO[11]  (.A(i[8]), .B(\cs[10]_net_1 ), .C(cs4), .Y(
        \cs_RNO_0[11] ));
    NOR2 \cs_RNO_1[3]  (.A(i[4]), .B(en1), .Y(N_236));
    OR2 en2_RNIA134 (.A(en2_net_1), .B(en1), .Y(sd_acq_en_c));
    NOR2 \cs_RNI1581[11]  (.A(ns_0_1_i_a2_1), .B(ns_0_1_i_a2_0), .Y(
        N_245));
    DFN1 \cs[12]  (.D(N_187_i_0), .CLK(ddsclkout_c), .Q(\cs[12]_net_1 )
        );
    VCC VCC_i (.Y(VCC));
    OR2 \cs_RNIGTQ[11]  (.A(\cs[4]_net_1 ), .B(\cs[11]_net_1 ), .Y(
        ns_0_1_i_a2_0));
    DFN1 \cs[3]  (.D(\cs_RNO_2[3] ), .CLK(ddsclkout_c), .Q(en1));
    NOR2A \cs_RNO[7]  (.A(cs4), .B(N_203), .Y(\cs_nsss[7] ));
    NOR2A \cs_RNO[1]  (.A(cs4), .B(\cs_i[0]_net_1 ), .Y(\cs_RNO_1[1] ));
    NOR2 \cs_RNO_1[8]  (.A(i[6]), .B(\cs[8]_net_1 ), .Y(N_222));
    OA1 \cs_RNO[9]  (.A(N_207), .B(\cs[9]_net_1 ), .C(
        \cs_srsts_0_i_0[9] ), .Y(N_182_i_0));
    DFN1 \cs[5]  (.D(\cs_RNO_2[5] ), .CLK(ddsclkout_c), .Q(
        \cs[5]_net_1 ));
    NOR2B cs4_0_o2 (.A(i_4[0]), .B(net_27), .Y(cs4));
    OR2 \cs_RNIH7D[14]  (.A(\cs[14]_net_1 ), .B(\cs[15]_net_1 ), .Y(
        ns_0_1_i_a2_1));
    OA1C \cs_RNO_0[3]  (.A(en1), .B(i[5]), .C(\cs[2]_net_1 ), .Y(N_237)
        );
    NOR3A \cs_RNO[8]  (.A(cs4), .B(N_221), .C(N_222), .Y(
        \cs_RNO_0[8]_net_1 ));
    DFN1 \cs[11]  (.D(\cs_RNO_0[11] ), .CLK(ddsclkout_c), .Q(
        \cs[11]_net_1 ));
    OA1A \cs_RNO_1[9]  (.A(i[7]), .B(\cs[5]_net_1 ), .C(cs4), .Y(
        \cs_srsts_0_i_0[9] ));
    DFN1 \cs[13]  (.D(\cs_nsss[13] ), .CLK(ddsclkout_c), .Q(
        \cs[13]_net_1 ));
    DFN1 \cs[2]  (.D(\cs_RNO_0[2]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[2]_net_1 ));
    NOR2B \cs_RNIRKL6[12]  (.A(i[9]), .B(\cs[12]_net_1 ), .Y(N_230));
    AOI1 \cs_RNO_0[8]  (.A(i_3[2]), .B(\cs[8]_net_1 ), .C(
        \cs[7]_net_1 ), .Y(N_221));
    OA1 \cs_RNO[12]  (.A(\cs_RNO_0[12]_net_1 ), .B(\cs[12]_net_1 ), .C(
        \cs_srsts_0_i_0[12] ), .Y(N_187_i_0));
    NOR2B \cs_RNITI37[6]  (.A(i[4]), .B(\cs[6]_net_1 ), .Y(N_234));
    NOR2A \cs_RNI4I52[13]  (.A(\cs[13]_net_1 ), .B(i[10]), .Y(N_231));
    AOI1B en2_RNO (.A(en2_0_0_o3_0), .B(N_203), .C(cs4), .Y(
        en2_RNO_net_1));
    GND GND_i (.Y(GND));
    NOR2 \cs_RNIV6R8[12]  (.A(N_231), .B(N_230), .Y(N_201));
    NOR3C \cs_RNO[14]  (.A(i[10]), .B(\cs[13]_net_1 ), .C(cs4), .Y(
        \cs_RNO[14]_net_1 ));
    DFN1 \cs[15]  (.D(\cs_RNO[15]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[15]_net_1 ));
    NOR2A \cs_RNO[15]  (.A(cs4), .B(N_245), .Y(\cs_RNO[15]_net_1 ));
    DFN1 \cs_i[0]  (.D(cs4), .CLK(ddsclkout_c), .Q(\cs_i[0]_net_1 ));
    DFN1 stateover (.D(stateover_RNO_0), .CLK(ddsclkout_c), .Q(
        sd_sacq_state_0_stateover));
    DFN1 \cs[10]  (.D(\cs_nsss[10] ), .CLK(ddsclkout_c), .Q(
        \cs[10]_net_1 ));
    NOR3A en2_RNO_0 (.A(N_201), .B(N_232), .C(N_233), .Y(en2_0_0_o3_0));
    AOI1 \cs_RNO_0[6]  (.A(i_3[2]), .B(\cs[5]_net_1 ), .C(
        \cs[6]_net_1 ), .Y(N_218));
    NOR3A \cs_RNO[2]  (.A(cs4), .B(N_214), .C(N_215), .Y(
        \cs_RNO_0[2]_net_1 ));
    OA1C \cs_RNO_0[2]  (.A(\cs[2]_net_1 ), .B(i[4]), .C(\cs[1]_net_1 ), 
        .Y(N_214));
    AO1B stateover_RNO (.A(sd_sacq_state_0_stateover), .B(N_245), .C(
        cs4), .Y(stateover_RNO_0));
    NOR3B \cs_RNO_0[12]  (.A(\cs[5]_net_1 ), .B(i_3[3]), .C(i_3[2]), 
        .Y(\cs_RNO_0[12]_net_1 ));
    NOR2A \cs_RNI0N37[7]  (.A(\cs[7]_net_1 ), .B(i[6]), .Y(N_235));
    NOR2 \cs_RNO_1[5]  (.A(i_4[1]), .B(\cs[8]_net_1 ), .Y(N_217));
    NOR3C \cs_RNO[4]  (.A(en1), .B(i[5]), .C(cs4), .Y(\cs_RNO_1[4] ));
    DFN1 \cs[9]  (.D(N_182_i_0), .CLK(ddsclkout_c), .Q(\cs[9]_net_1 ));
    OA1C \cs_RNO_0[5]  (.A(\cs[8]_net_1 ), .B(i_3[2]), .C(
        \cs[1]_net_1 ), .Y(N_216));
    DFN1 \cs[8]  (.D(\cs_RNO_0[8]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[8]_net_1 ));
    NOR2A \cs_RNO_1[6]  (.A(i[4]), .B(\cs[5]_net_1 ), .Y(N_219));
    NOR3A \cs_RNO[6]  (.A(cs4), .B(N_218), .C(N_219), .Y(
        \cs_RNO_1[6]_net_1 ));
    NOR2A \cs_RNO_1[2]  (.A(i_4[1]), .B(\cs[2]_net_1 ), .Y(N_215));
    NOR2A \cs_RNIOKL6[10]  (.A(\cs[10]_net_1 ), .B(i[8]), .Y(N_233));
    DFN1 \cs[14]  (.D(\cs_RNO[14]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[14]_net_1 ));
    NOR3A \cs_RNO[3]  (.A(cs4), .B(N_237), .C(N_236), .Y(\cs_RNO_2[3] )
        );
    DFN1 \cs[1]  (.D(\cs_RNO_1[1] ), .CLK(ddsclkout_c), .Q(
        \cs[1]_net_1 ));
    OA1A \cs_RNO_1[12]  (.A(i[9]), .B(\cs[5]_net_1 ), .C(cs4), .Y(
        \cs_srsts_0_i_0[12] ));
    NOR3A \cs_RNO[5]  (.A(cs4), .B(N_216), .C(N_217), .Y(\cs_RNO_2[5] )
        );
    DFN1 \cs[4]  (.D(\cs_RNO_1[4] ), .CLK(ddsclkout_c), .Q(
        \cs[4]_net_1 ));
    DFN1 \cs[7]  (.D(\cs_nsss[7] ), .CLK(ddsclkout_c), .Q(
        \cs[7]_net_1 ));
    DFN1 en2 (.D(en2_RNO_net_1), .CLK(ddsclkout_c), .Q(en2_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR3A \cs_RNO_0[9]  (.A(\cs[5]_net_1 ), .B(i_3[2]), .C(i_3[3]), .Y(
        N_207));
    
endmodule


module sd_sacq_inc(
       count_1,
       count,
       count_4,
       count1
    );
input  [7:5] count_1;
input  [21:8] count;
input  [4:0] count_4;
output [21:1] count1;

    wire Rcout_4_net, Rcout_6_net, inc_2_net, inc_5_net, Rcout_16_net, 
        Rcout_5_net, inc_8_net, inc_1_net, Rcout_8_net, Rcout_7_net, 
        Rcout_17_net, inc_17_net, inc1_25_net, inc_16_net, 
        Rcout_18_net, incb_17_net, inc_28_net, incb_16_net, inc_22_net, 
        inc_27_net, Rcout_19_net, Rcout_9_net, incb_2_net, inc_10_net, 
        incb_5_net, inc_12_net, Rcout_13_net, Rcout_10_net, 
        Rcout_15_net, Rcout_11_net, inc_14_net, Rcout_12_net, 
        Rcout_14_net, inc_20_net, inc_24_net, Rcout_20_net, inc_31_net, 
        Rcout_21_net, inc_33_net, GND, VCC, GND_0, VCC_0;
    
    AND3 QAND2_26_inst (.A(incb_17_net), .B(inc_28_net), .C(inc_31_net)
        , .Y(Rcout_20_net));
    AND3 AND2b_9_inst (.A(count_4[0]), .B(count_4[1]), .C(count_4[2]), 
        .Y(incb_2_net));
    AND3 FND2_9_inst (.A(inc_12_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_10_net));
    AND2 AND2_4_inst (.A(inc_2_net), .B(count_4[3]), .Y(Rcout_4_net));
    XOR2 YXOR2_14_inst (.A(Rcout_18_net), .B(count[18]), .Y(count1[18])
        );
    AND3 PAND2_19_inst (.A(inc_22_net), .B(inc_16_net), .C(count[16]), 
        .Y(inc1_25_net));
    AND3 AND2_15_inst (.A(inc_16_net), .B(inc_17_net), .C(inc_20_net), 
        .Y(Rcout_14_net));
    AND3 AND2_1_12_inst (.A(incb_2_net), .B(incb_5_net), .C(inc_10_net)
        , .Y(inc_17_net));
    AND2 AND2_13_inst (.A(inc_17_net), .B(inc_16_net), .Y(Rcout_12_net)
        );
    AND3 VAND2_18_inst (.A(inc_17_net), .B(inc_24_net), .C(count[15]), 
        .Y(Rcout_16_net));
    AND3 AND2_12_inst (.A(count[9]), .B(count[10]), .C(count[11]), .Y(
        inc_16_net));
    AND2 VAND2_17_inst (.A(inc_22_net), .B(inc_16_net), .Y(inc_24_net));
    XOR2 QXOR2_16_inst (.A(Rcout_20_net), .B(count[20]), .Y(count1[20])
        );
    AND2 YAND2_23_inst (.A(incb_17_net), .B(inc_28_net), .Y(
        Rcout_18_net));
    VCC VCC_i (.Y(VCC));
    AND3 AND2_1_7_inst (.A(inc_2_net), .B(inc_5_net), .C(count_1[6]), 
        .Y(Rcout_7_net));
    XOR2 HOR2_10_inst (.A(Rcout_13_net), .B(count[13]), .Y(count1[13]));
    AND3 AND2_1_8_inst (.A(inc_2_net), .B(inc_5_net), .C(inc_8_net), 
        .Y(Rcout_8_net));
    XOR2 XOR2_4_inst (.A(Rcout_5_net), .B(count_1[5]), .Y(count1[5]));
    XOR2 SXOR2_17_inst (.A(Rcout_21_net), .B(count[21]), .Y(count1[21])
        );
    AND3 SAND2_28_inst (.A(incb_17_net), .B(inc_28_net), .C(inc_33_net)
        , .Y(Rcout_21_net));
    AND3 SAND2_27_inst (.A(count[18]), .B(count[19]), .C(count[20]), 
        .Y(inc_33_net));
    AND3 OAND2_24_inst (.A(incb_17_net), .B(inc_28_net), .C(count[18]), 
        .Y(Rcout_19_net));
    AND2 AND2_7_inst (.A(inc_2_net), .B(inc_5_net), .Y(Rcout_6_net));
    AND2 AND2_14_inst (.A(count[12]), .B(count[13]), .Y(inc_20_net));
    XOR2 VXOR2_13_inst (.A(Rcout_16_net), .B(count[16]), .Y(count1[16])
        );
    AND3 TND2_15_inst (.A(inc_16_net), .B(inc_17_net), .C(inc_22_net), 
        .Y(Rcout_15_net));
    XOR2 XOR2_3_inst (.A(Rcout_4_net), .B(count_4[4]), .Y(count1[4]));
    AND2 FND2_8_inst (.A(incb_2_net), .B(count[9]), .Y(inc_12_net));
    XOR2 XOR2_7_inst (.A(Rcout_9_net), .B(count[9]), .Y(count1[9]));
    XOR2 UXOR2_12_inst (.A(Rcout_15_net), .B(count[15]), .Y(count1[15])
        );
    AND3 AND2_9_inst (.A(count_1[6]), .B(count_1[7]), .C(count[8]), .Y(
        inc_10_net));
    GND GND_i (.Y(GND));
    AND3 AND2_11_inst (.A(inc_14_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_11_net));
    XOR2 XOR2_6_inst (.A(Rcout_8_net), .B(count[8]), .Y(count1[8]));
    AND3 YAND2B_22_inst (.A(incb_2_net), .B(incb_5_net), .C(inc_10_net)
        , .Y(incb_17_net));
    XOR2 XOR2_1_5_inst (.A(Rcout_7_net), .B(count_1[7]), .Y(count1[7]));
    AND2 QAND2_25_inst (.A(count[18]), .B(count[19]), .Y(inc_31_net));
    AND3 TAND2_15_inst (.A(count[12]), .B(count[13]), .C(count[14]), 
        .Y(inc_22_net));
    AND3 AND2_3_inst (.A(count_4[0]), .B(count_4[1]), .C(count_4[2]), 
        .Y(inc_2_net));
    AND3 YAND2_22_inst (.A(incb_16_net), .B(inc_22_net), .C(inc_27_net)
        , .Y(inc_28_net));
    AND3 fAND2_8_inst (.A(incb_2_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_9_net));
    AND3 AND2_6_inst (.A(count_4[3]), .B(count_4[4]), .C(count_1[5]), 
        .Y(inc_5_net));
    AND3 AND2b_12_inst (.A(count_4[3]), .B(count_4[4]), .C(count_1[5]), 
        .Y(incb_5_net));
    XOR2 XOR2_2_1_inst (.A(inc_1_net), .B(count_4[2]), .Y(count1[2]));
    AND3 YAND2BB_21_inst (.A(count[9]), .B(count[10]), .C(count[11]), 
        .Y(incb_16_net));
    XOR2 XOR2_1_inst (.A(count_4[0]), .B(count_4[1]), .Y(count1[1]));
    XOR2 OXOR2_15_inst (.A(Rcout_19_net), .B(count[19]), .Y(count1[19])
        );
    XOR2 XOR2_9_inst (.A(Rcout_11_net), .B(count[11]), .Y(count1[11]));
    XOR2 PXOR2_13_inst (.A(Rcout_17_net), .B(count[17]), .Y(count1[17])
        );
    AND3 YAND2_21_inst (.A(count[15]), .B(count[16]), .C(count[17]), 
        .Y(inc_27_net));
    XOR2 XOR2_2_inst (.A(inc_2_net), .B(count_4[3]), .Y(count1[3]));
    AND3 PAND2_20_inst (.A(inc_17_net), .B(inc1_25_net), .C(count[15]), 
        .Y(Rcout_17_net));
    AND2 AND2_8_inst (.A(count_1[6]), .B(count_1[7]), .Y(inc_8_net));
    AND3 HND2_13_inst (.A(inc_17_net), .B(inc_16_net), .C(count[12]), 
        .Y(Rcout_13_net));
    XOR2 POR2_9_inst (.A(Rcout_12_net), .B(count[12]), .Y(count1[12]));
    XOR2 XOR2_5_inst (.A(Rcout_6_net), .B(count_1[6]), .Y(count1[6]));
    AND2 AND2_2_inst (.A(count_4[0]), .B(count_4[1]), .Y(inc_1_net));
    AND3 AND2_5_inst (.A(inc_2_net), .B(count_4[3]), .C(count_4[4]), 
        .Y(Rcout_5_net));
    XOR2 FOR2_8_inst (.A(Rcout_10_net), .B(count[10]), .Y(count1[10]));
    XOR2 XOR2_11_inst (.A(Rcout_14_net), .B(count[14]), .Y(count1[14]));
    AND3 AND2_10_inst (.A(incb_2_net), .B(count[9]), .C(count[10]), .Y(
        inc_14_net));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module sd_sacq_timer(
       count,
       count_1,
       count_4,
       net_27,
       ddsclkout_c,
       sd_sacq_state_0_stateover,
       scalestate_0_s_acq
    );
output [21:8] count;
output [7:5] count_1;
output [4:0] count_4;
input  net_27;
input  ddsclkout_c;
input  sd_sacq_state_0_stateover;
input  scalestate_0_s_acq;

    wire \count_3[0] , \count_3[1] , \count1[1] , \count_3[2] , 
        \count1[2] , \count_3[3] , \count1[3] , \count_3[4] , 
        \count1[4] , \count_3[5] , \count1[5] , \count_3[6] , 
        \count1[6] , \count_3[7] , \count1[7] , \count_3[8] , 
        \count1[8] , \count_3[9] , \count1[9] , \count_3[10] , 
        \count1[10] , \count_3[11] , \count1[11] , \count_3[12] , 
        \count1[12] , \count_3[13] , \count1[13] , \count_3[14] , 
        \count1[14] , \count_3[15] , \count1[15] , \count_3[16] , 
        \count1[16] , \count_3[17] , \count1[17] , \count_3[18] , 
        \count1[18] , \count_3[19] , \count1[19] , \count_3[20] , 
        \count1[20] , \count_3[21] , \count1[21] , GND, VCC, GND_0, 
        VCC_0;
    
    NOR3C \count_RNO[21]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[21] ), .Y(\count_3[21] )
        );
    DFN1C0 \count[5]  (.D(\count_3[5] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_1[5]));
    DFN1C0 \count[1]  (.D(\count_3[1] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_4[1]));
    DFN1C0 \count[10]  (.D(\count_3[10] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[10]));
    DFN1C0 \count[0]  (.D(\count_3[0] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_4[0]));
    DFN1C0 \count[14]  (.D(\count_3[14] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[14]));
    NOR3C \count_RNO[7]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[7] ), .Y(\count_3[7] ));
    NOR3C \count_RNO[15]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[15] ), .Y(\count_3[15] )
        );
    NOR3C \count_RNO[2]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[2] ), .Y(\count_3[2] ));
    NOR3C \count_RNO[9]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[9] ), .Y(\count_3[9] ));
    DFN1C0 \count[20]  (.D(\count_3[20] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[20]));
    VCC VCC_i (.Y(VCC));
    NOR3C \count_RNO[4]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[4] ), .Y(\count_3[4] ));
    DFN1C0 \count[8]  (.D(\count_3[8] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[8]));
    NOR3C \count_RNO[10]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[10] ), .Y(\count_3[10] )
        );
    DFN1C0 \count[19]  (.D(\count_3[19] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[19]));
    DFN1C0 \count[15]  (.D(\count_3[15] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[15]));
    NOR3C \count_RNO[3]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[3] ), .Y(\count_3[3] ));
    DFN1C0 \count[11]  (.D(\count_3[11] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[11]));
    sd_sacq_inc sd_sacq_inc_0 (.count_1({count_1[7], count_1[6], 
        count_1[5]}), .count({count[21], count[20], count[19], 
        count[18], count[17], count[16], count[15], count[14], 
        count[13], count[12], count[11], count[10], count[9], count[8]})
        , .count_4({count_4[4], count_4[3], count_4[2], count_4[1], 
        count_4[0]}), .count1({\count1[21] , \count1[20] , 
        \count1[19] , \count1[18] , \count1[17] , \count1[16] , 
        \count1[15] , \count1[14] , \count1[13] , \count1[12] , 
        \count1[11] , \count1[10] , \count1[9] , \count1[8] , 
        \count1[7] , \count1[6] , \count1[5] , \count1[4] , 
        \count1[3] , \count1[2] , \count1[1] }));
    NOR3C \count_RNO[8]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[8] ), .Y(\count_3[8] ));
    DFN1C0 \count[13]  (.D(\count_3[13] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[13]));
    NOR3C \count_RNO[5]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[5] ), .Y(\count_3[5] ));
    NOR3C \count_RNO[1]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[1] ), .Y(\count_3[1] ));
    NOR3C \count_RNO[11]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[11] ), .Y(\count_3[11] )
        );
    DFN1C0 \count[2]  (.D(\count_3[2] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_4[2]));
    DFN1C0 \count[21]  (.D(\count_3[21] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[21]));
    NOR3C \count_RNO[16]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[16] ), .Y(\count_3[16] )
        );
    GND GND_i (.Y(GND));
    DFN1C0 \count[9]  (.D(\count_3[9] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[9]));
    DFN1C0 \count[16]  (.D(\count_3[16] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[16]));
    NOR3C \count_RNO[6]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[6] ), .Y(\count_3[6] ));
    NOR3C \count_RNO[12]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[12] ), .Y(\count_3[12] )
        );
    NOR3B \count_RNO[0]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(count_4[0]), .Y(\count_3[0] ));
    DFN1C0 \count[6]  (.D(\count_3[6] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_1[6]));
    DFN1C0 \count[3]  (.D(\count_3[3] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_4[3]));
    NOR3C \count_RNO[17]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[17] ), .Y(\count_3[17] )
        );
    NOR3C \count_RNO[14]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[14] ), .Y(\count_3[14] )
        );
    NOR3C \count_RNO[19]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[19] ), .Y(\count_3[19] )
        );
    NOR3C \count_RNO[18]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[18] ), .Y(\count_3[18] )
        );
    NOR3C \count_RNO[13]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[13] ), .Y(\count_3[13] )
        );
    DFN1C0 \count[18]  (.D(\count_3[18] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[18]));
    NOR3C \count_RNO[20]  (.A(scalestate_0_s_acq), .B(
        sd_sacq_state_0_stateover), .C(\count1[20] ), .Y(\count_3[20] )
        );
    DFN1C0 \count[17]  (.D(\count_3[17] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[17]));
    DFN1C0 \count[4]  (.D(\count_3[4] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_4[4]));
    DFN1C0 \count[12]  (.D(\count_3[12] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count[12]));
    DFN1C0 \count[7]  (.D(\count_3[7] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_1[7]));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module sd_acq_top(
       sd_sacq_choice,
       sd_sacq_data,
       i_4_1,
       i_0_0,
       sd_acq_en_c,
       net_27,
       scalestate_0_s_acq,
       top_code_0_sd_sacq_load,
       s_acq180_c,
       scalestate_0_long_opentime,
       GLA,
       ddsclkout_c
    );
input  [3:0] sd_sacq_choice;
input  [15:0] sd_sacq_data;
output i_4_1;
input  [1:1] i_0_0;
output sd_acq_en_c;
input  net_27;
input  scalestate_0_s_acq;
input  top_code_0_sd_sacq_load;
input  s_acq180_c;
input  scalestate_0_long_opentime;
input  GLA;
input  ddsclkout_c;

    wire \i[4] , \i[5] , \i[6] , \i[7] , \i[8] , \i[9] , \i[10] , 
        \i_3[2] , \i_3[3] , \i_4[0] , \count_4[0] , \count_4[1] , 
        \count_4[2] , \count_4[3] , \count_4[4] , \count_1[5] , 
        \count_1[6] , \count_1[7] , \count[8] , \count[9] , 
        \count[10] , \count[11] , \count[12] , \count[13] , 
        \count[14] , \count[15] , \count[16] , \count[17] , 
        \count[18] , \count[19] , \count[20] , \count[21] , 
        sd_sacq_state_0_stateover, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    sd_sacq_coder sd_sacq_coder_0 (.i({\i[10] , \i[9] , \i[8] , \i[7] , 
        \i[6] , \i[5] , \i[4] }), .i_3({\i_3[3] , \i_3[2] }), .i_0_0_0(
        i_0_0[1]), .i_4({i_4_1, \i_4[0] }), .sd_sacq_data({
        sd_sacq_data[15], sd_sacq_data[14], sd_sacq_data[13], 
        sd_sacq_data[12], sd_sacq_data[11], sd_sacq_data[10], 
        sd_sacq_data[9], sd_sacq_data[8], sd_sacq_data[7], 
        sd_sacq_data[6], sd_sacq_data[5], sd_sacq_data[4], 
        sd_sacq_data[3], sd_sacq_data[2], sd_sacq_data[1], 
        sd_sacq_data[0]}), .sd_sacq_choice({sd_sacq_choice[3], 
        sd_sacq_choice[2], sd_sacq_choice[1], sd_sacq_choice[0]}), 
        .count_4({\count_4[4] , \count_4[3] , \count_4[2] , 
        \count_4[1] , \count_4[0] }), .count_1({\count_1[7] , 
        \count_1[6] , \count_1[5] }), .count({\count[21] , \count[20] , 
        \count[19] , \count[18] , \count[17] , \count[16] , 
        \count[15] , \count[14] , \count[13] , \count[12] , 
        \count[11] , \count[10] , \count[9] , \count[8] }), 
        .ddsclkout_c(ddsclkout_c), .GLA(GLA), 
        .scalestate_0_long_opentime(scalestate_0_long_opentime), 
        .s_acq180_c(s_acq180_c), .top_code_0_sd_sacq_load(
        top_code_0_sd_sacq_load), .scalestate_0_s_acq(
        scalestate_0_s_acq), .net_27(net_27));
    sd_sacq_state sd_sacq_state_0 (.i_3({\i_3[3] , \i_3[2] }), .i_4({
        i_4_1, \i_4[0] }), .i({\i[10] , \i[9] , \i[8] , \i[7] , \i[6] , 
        \i[5] , \i[4] }), .ddsclkout_c(ddsclkout_c), .sd_acq_en_c(
        sd_acq_en_c), .sd_sacq_state_0_stateover(
        sd_sacq_state_0_stateover), .net_27(net_27));
    GND GND_i_0 (.Y(GND_0));
    sd_sacq_timer sd_sacq_timer_0 (.count({\count[21] , \count[20] , 
        \count[19] , \count[18] , \count[17] , \count[16] , 
        \count[15] , \count[14] , \count[13] , \count[12] , 
        \count[11] , \count[10] , \count[9] , \count[8] }), .count_1({
        \count_1[7] , \count_1[6] , \count_1[5] }), .count_4({
        \count_4[4] , \count_4[3] , \count_4[2] , \count_4[1] , 
        \count_4[0] }), .net_27(net_27), .ddsclkout_c(ddsclkout_c), 
        .sd_sacq_state_0_stateover(sd_sacq_state_0_stateover), 
        .scalestate_0_s_acq(scalestate_0_s_acq));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_2(
       un1_off_on_coder_0,
       GLA,
       DUMP_OFF_1_dump_off,
       off_on_state_0_state_over,
       nsctrl_choice_0_dumponoff_rst
    );
input  [1:0] un1_off_on_coder_0;
input  GLA;
output DUMP_OFF_1_dump_off;
output off_on_state_0_state_over;
input  nsctrl_choice_0_dumponoff_rst;

    wire state_over_1_0, N_14, N_42, \cs_nsss[0] , \cs_nsss[1] , 
        \cs_ns[1] , \cs[1]_net_1 , GND, VCC, GND_0, VCC_0;
    
    NOR2B state_over_RNO_0 (.A(un1_off_on_coder_0[0]), .B(
        nsctrl_choice_0_dumponoff_rst), .Y(state_over_1_0));
    DFN1 state_over (.D(N_14), .CLK(GLA), .Q(off_on_state_0_state_over)
        );
    AOI1 \cs_RNILT8E[1]  (.A(DUMP_OFF_1_dump_off), .B(
        un1_off_on_coder_0[1]), .C(\cs[1]_net_1 ), .Y(N_42));
    DFN1 \cs[0]  (.D(\cs_nsss[0] ), .CLK(GLA), .Q(DUMP_OFF_1_dump_off));
    NOR3C \cs_RNO[0]  (.A(N_42), .B(nsctrl_choice_0_dumponoff_rst), .C(
        un1_off_on_coder_0[0]), .Y(\cs_nsss[0] ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 \cs[1]  (.D(\cs_nsss[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3C \cs_RNO[1]  (.A(\cs_ns[1] ), .B(
        nsctrl_choice_0_dumponoff_rst), .C(un1_off_on_coder_0[0]), .Y(
        \cs_nsss[1] ));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    MX2 \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(un1_off_on_coder_0[1]), 
        .S(DUMP_OFF_1_dump_off), .Y(\cs_ns[1] ));
    AO1B state_over_RNO (.A(off_on_state_0_state_over), .B(N_42), .C(
        state_over_1_0), .Y(N_14));
    
endmodule


module off_on_coder_2(
       un1_off_on_coder_0,
       un1_off_on_timer_0,
       GLA,
       nsctrl_choice_0_dumpoff_ctr,
       nsctrl_choice_0_dumponoff_rst
    );
output [1:0] un1_off_on_coder_0;
input  [4:0] un1_off_on_timer_0;
input  GLA;
input  nsctrl_choice_0_dumpoff_ctr;
input  nsctrl_choice_0_dumponoff_rst;

    wire \i_0_1[1] , N_4, N_17, N_3, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    NOR3B \i_RNO_1[1]  (.A(un1_off_on_timer_0[2]), .B(
        un1_off_on_timer_0[4]), .C(un1_off_on_timer_0[3]), .Y(
        \i_0_1[1] ));
    DFN1 \i[1]  (.D(N_4), .CLK(GLA), .Q(un1_off_on_coder_0[1]));
    GND GND_i_0 (.Y(GND_0));
    NOR3C \i_RNO[1]  (.A(nsctrl_choice_0_dumponoff_rst), .B(N_17), .C(
        \i_0_1[1] ), .Y(N_4));
    VCC VCC_i (.Y(VCC));
    NOR2 \i_RNO_0[1]  (.A(un1_off_on_timer_0[1]), .B(
        un1_off_on_timer_0[0]), .Y(N_17));
    NOR2B \i_RNO[0]  (.A(nsctrl_choice_0_dumponoff_rst), .B(
        nsctrl_choice_0_dumpoff_ctr), .Y(N_3));
    DFN1 \i[0]  (.D(N_3), .CLK(GLA), .Q(un1_off_on_coder_0[0]));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_2(
       un1_off_on_timer_0,
       GLA,
       nsctrl_choice_0_dumponoff_rst,
       off_on_state_0_state_over,
       nsctrl_choice_0_dumpoff_ctr
    );
output [4:0] un1_off_on_timer_0;
input  GLA;
input  nsctrl_choice_0_dumponoff_rst;
input  off_on_state_0_state_over;
input  nsctrl_choice_0_dumpoff_ctr;

    wire count_0_sqmuxa_net_1, N_9, N_13, N_7, N_12, N_5, N_15_i, N_11, 
        count_n0, GND, VCC, GND_0, VCC_0;
    
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(un1_off_on_timer_0[0]), .B(
        un1_off_on_timer_0[1]), .C(count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(un1_off_on_timer_0[3]));
    NOR2B \count_RNIB785[1]  (.A(un1_off_on_timer_0[1]), .B(
        un1_off_on_timer_0[0]), .Y(N_12));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(un1_off_on_timer_0[0])
        );
    XA1B \count_RNO[3]  (.A(N_13), .B(un1_off_on_timer_0[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    AX1E \count_RNO_0[4]  (.A(N_13), .B(un1_off_on_timer_0[3]), .C(
        un1_off_on_timer_0[4]), .Y(N_15_i));
    XA1B \count_RNO[2]  (.A(N_12), .B(un1_off_on_timer_0[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(nsctrl_choice_0_dumpoff_ctr), .B(
        off_on_state_0_state_over), .C(nsctrl_choice_0_dumponoff_rst), 
        .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \count_RNO[4]  (.A(count_0_sqmuxa_net_1), .B(N_15_i), .Y(N_11)
        );
    NOR2B \count_RNI2HS7[2]  (.A(un1_off_on_timer_0[2]), .B(N_12), .Y(
        N_13));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(un1_off_on_timer_0[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(un1_off_on_timer_0[4]));
    NOR2 \count_RNO[0]  (.A(un1_off_on_timer_0[0]), .B(
        count_0_sqmuxa_net_1), .Y(count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(un1_off_on_timer_0[2]));
    
endmodule


module DUMP_OFF_DUMP_OFF_0_1(
       nsctrl_choice_0_dumpoff_ctr,
       nsctrl_choice_0_dumponoff_rst,
       DUMP_OFF_1_dump_off,
       GLA
    );
input  nsctrl_choice_0_dumpoff_ctr;
input  nsctrl_choice_0_dumponoff_rst;
output DUMP_OFF_1_dump_off;
input  GLA;

    wire \un1_off_on_coder_0[0] , \un1_off_on_coder_0[1] , 
        off_on_state_0_state_over, \un1_off_on_timer_0[0] , 
        \un1_off_on_timer_0[1] , \un1_off_on_timer_0[2] , 
        \un1_off_on_timer_0[3] , \un1_off_on_timer_0[4] , GND, VCC, 
        GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_2 
        off_on_state_0 (.un1_off_on_coder_0({\un1_off_on_coder_0[1] , 
        \un1_off_on_coder_0[0] }), .GLA(GLA), .DUMP_OFF_1_dump_off(
        DUMP_OFF_1_dump_off), .off_on_state_0_state_over(
        off_on_state_0_state_over), .nsctrl_choice_0_dumponoff_rst(
        nsctrl_choice_0_dumponoff_rst));
    off_on_coder_2 off_on_coder_0 (.un1_off_on_coder_0({
        \un1_off_on_coder_0[1] , \un1_off_on_coder_0[0] }), 
        .un1_off_on_timer_0({\un1_off_on_timer_0[4] , 
        \un1_off_on_timer_0[3] , \un1_off_on_timer_0[2] , 
        \un1_off_on_timer_0[1] , \un1_off_on_timer_0[0] }), .GLA(GLA), 
        .nsctrl_choice_0_dumpoff_ctr(nsctrl_choice_0_dumpoff_ctr), 
        .nsctrl_choice_0_dumponoff_rst(nsctrl_choice_0_dumponoff_rst));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_2 
        off_on_timer_0 (.un1_off_on_timer_0({\un1_off_on_timer_0[4] , 
        \un1_off_on_timer_0[3] , \un1_off_on_timer_0[2] , 
        \un1_off_on_timer_0[1] , \un1_off_on_timer_0[0] }), .GLA(GLA), 
        .nsctrl_choice_0_dumponoff_rst(nsctrl_choice_0_dumponoff_rst), 
        .off_on_state_0_state_over(off_on_state_0_state_over), 
        .nsctrl_choice_0_dumpoff_ctr(nsctrl_choice_0_dumpoff_ctr));
    GND GND_i (.Y(GND));
    
endmodule


module necount_cmp(
       M_NUM,
       necount,
       necount_LE_M_1
    );
input  [11:0] M_NUM;
input  [11:0] necount;
output necount_LE_M_1;

    wire AND3_3_Y, XNOR2_2_Y, XNOR2_1_Y, XNOR2_10_Y, OR2A_7_Y, 
        NAND3A_4_Y, OR2A_1_Y, NAND3A_7_Y, OR2A_2_Y, OR2A_4_Y, 
        XNOR2_6_Y, XNOR2_7_Y, AO1_0_Y, NAND3A_1_Y, NAND3A_6_Y, 
        NAND3A_0_Y, NOR3A_0_Y, NAND3A_2_Y, XNOR2_0_Y, OR2A_6_Y, 
        NOR3A_1_Y, AO1C_1_Y, OR2A_3_Y, XNOR2_9_Y, AO1_1_Y, AND3_2_Y, 
        NAND3A_5_Y, XNOR2_4_Y, NOR3A_2_Y, NAND3A_3_Y, XNOR2_8_Y, 
        AND3_1_Y, XNOR2_5_Y, XNOR2_3_Y, OR2A_0_Y, NOR3A_3_Y, AND3_0_Y, 
        AND2_0_Y, OR2A_5_Y, AO1C_0_Y, XNOR2_11_Y, AO1C_2_Y, AO1C_3_Y, 
        GND, VCC, GND_0, VCC_0;
    
    OR2A OR2A_1 (.A(M_NUM[11]), .B(necount[11]), .Y(OR2A_1_Y));
    XNOR2 XNOR2_3 (.A(necount[8]), .B(M_NUM[8]), .Y(XNOR2_3_Y));
    NAND3A NAND3A_2 (.A(M_NUM[4]), .B(necount[4]), .C(OR2A_0_Y), .Y(
        NAND3A_2_Y));
    NAND3A NAND3A_6 (.A(NOR3A_1_Y), .B(OR2A_6_Y), .C(NAND3A_4_Y), .Y(
        NAND3A_6_Y));
    NOR3A NOR3A_1 (.A(OR2A_1_Y), .B(AO1C_0_Y), .C(M_NUM[9]), .Y(
        NOR3A_1_Y));
    AND3 AND3_2 (.A(XNOR2_0_Y), .B(XNOR2_11_Y), .C(XNOR2_8_Y), .Y(
        AND3_2_Y));
    AO1C AO1C_3 (.A(necount[4]), .B(M_NUM[4]), .C(necount[3]), .Y(
        AO1C_3_Y));
    AND2 AND2_0 (.A(XNOR2_4_Y), .B(XNOR2_6_Y), .Y(AND2_0_Y));
    NOR3A NOR3A_2 (.A(OR2A_3_Y), .B(AO1C_2_Y), .C(M_NUM[6]), .Y(
        NOR3A_2_Y));
    VCC VCC_i (.Y(VCC));
    AO1 AO1_1 (.A(AND3_2_Y), .B(NAND3A_5_Y), .C(NAND3A_0_Y), .Y(
        AO1_1_Y));
    NAND3A NAND3A_4 (.A(M_NUM[10]), .B(necount[10]), .C(OR2A_1_Y), .Y(
        NAND3A_4_Y));
    XNOR2 XNOR2_9 (.A(necount[6]), .B(M_NUM[6]), .Y(XNOR2_9_Y));
    NAND3A NAND3A_1 (.A(NOR3A_2_Y), .B(OR2A_4_Y), .C(NAND3A_3_Y), .Y(
        NAND3A_1_Y));
    AND3 AND3_0 (.A(XNOR2_7_Y), .B(AND3_1_Y), .C(AND2_0_Y), .Y(
        AND3_0_Y));
    OR2A OR2A_3 (.A(M_NUM[8]), .B(necount[8]), .Y(OR2A_3_Y));
    XNOR2 XNOR2_4 (.A(necount[10]), .B(M_NUM[10]), .Y(XNOR2_4_Y));
    OR2A OR2A_6 (.A(necount[11]), .B(M_NUM[11]), .Y(OR2A_6_Y));
    AO1C AO1C_0 (.A(necount[10]), .B(M_NUM[10]), .C(necount[9]), .Y(
        AO1C_0_Y));
    XNOR2 XNOR2_1 (.A(M_NUM[10]), .B(necount[10]), .Y(XNOR2_1_Y));
    XNOR2 XNOR2_8 (.A(M_NUM[5]), .B(necount[5]), .Y(XNOR2_8_Y));
    XNOR2 XNOR2_5 (.A(necount[7]), .B(M_NUM[7]), .Y(XNOR2_5_Y));
    OR2A OR2A_7 (.A(necount[5]), .B(M_NUM[5]), .Y(OR2A_7_Y));
    XNOR2 XNOR2_6 (.A(necount[11]), .B(M_NUM[11]), .Y(XNOR2_6_Y));
    GND GND_i (.Y(GND));
    XNOR2 XNOR2_10 (.A(M_NUM[11]), .B(necount[11]), .Y(XNOR2_10_Y));
    NOR3A NOR3A_0 (.A(OR2A_0_Y), .B(AO1C_3_Y), .C(M_NUM[3]), .Y(
        NOR3A_0_Y));
    NAND3A NAND3A_3 (.A(M_NUM[7]), .B(necount[7]), .C(OR2A_3_Y), .Y(
        NAND3A_3_Y));
    XNOR2 XNOR2_2 (.A(M_NUM[9]), .B(necount[9]), .Y(XNOR2_2_Y));
    NAND3A NAND3A_5 (.A(NOR3A_3_Y), .B(OR2A_5_Y), .C(NAND3A_7_Y), .Y(
        NAND3A_5_Y));
    AND3 AND3_3 (.A(XNOR2_2_Y), .B(XNOR2_1_Y), .C(XNOR2_10_Y), .Y(
        AND3_3_Y));
    AND3 AND3_1 (.A(XNOR2_9_Y), .B(XNOR2_5_Y), .C(XNOR2_3_Y), .Y(
        AND3_1_Y));
    NAND3A NAND3A_7 (.A(M_NUM[1]), .B(necount[1]), .C(OR2A_2_Y), .Y(
        NAND3A_7_Y));
    OR2A OR2A_4 (.A(necount[8]), .B(M_NUM[8]), .Y(OR2A_4_Y));
    OR2A OR2A_0 (.A(M_NUM[5]), .B(necount[5]), .Y(OR2A_0_Y));
    AO1C AO1C_1 (.A(necount[1]), .B(M_NUM[1]), .C(necount[0]), .Y(
        AO1C_1_Y));
    XNOR2 XNOR2_11 (.A(M_NUM[4]), .B(necount[4]), .Y(XNOR2_11_Y));
    XNOR2 XNOR2_0 (.A(M_NUM[3]), .B(necount[3]), .Y(XNOR2_0_Y));
    OR2A OR2A_2 (.A(M_NUM[2]), .B(necount[2]), .Y(OR2A_2_Y));
    AO1C AO1C_2 (.A(necount[7]), .B(M_NUM[7]), .C(necount[6]), .Y(
        AO1C_2_Y));
    OR2A OR2A_5 (.A(necount[2]), .B(M_NUM[2]), .Y(OR2A_5_Y));
    AO1 AO1_0 (.A(AND3_3_Y), .B(NAND3A_1_Y), .C(NAND3A_6_Y), .Y(
        AO1_0_Y));
    NOR3A NOR3A_3 (.A(OR2A_2_Y), .B(AO1C_1_Y), .C(M_NUM[0]), .Y(
        NOR3A_3_Y));
    XNOR2 XNOR2_7 (.A(necount[9]), .B(M_NUM[9]), .Y(XNOR2_7_Y));
    NAND3A NAND3A_0 (.A(NOR3A_0_Y), .B(OR2A_7_Y), .C(NAND3A_2_Y), .Y(
        NAND3A_0_Y));
    AOI1 AOI1_ALEB (.A(AND3_0_Y), .B(AO1_1_Y), .C(AO1_0_Y), .Y(
        necount_LE_M_1));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module necount_inc(
       necount,
       necount1
    );
input  [11:0] necount;
output [11:1] necount1;

    wire Rcout_8_net, Rcout_5_net, inc_2_net, Rcout_6_net, inc_5_net, 
        Rcout_4_net, Rcout_10_net, inc_12_net, inc_10_net, Rcout_9_net, 
        incb_2_net, Rcout_11_net, inc_14_net, inc_1_net, inc_8_net, 
        Rcout_7_net, GND, VCC, GND_0, VCC_0;
    
    AND3 AND2b_9_inst (.A(necount[0]), .B(necount[1]), .C(necount[2]), 
        .Y(incb_2_net));
    AND3 AND2_5_inst (.A(inc_2_net), .B(necount[3]), .C(necount[4]), 
        .Y(Rcout_5_net));
    XOR2 XOR2_4_inst (.A(Rcout_5_net), .B(necount[5]), .Y(necount1[5]));
    XOR2 XOR2_1_inst (.A(necount[0]), .B(necount[1]), .Y(necount1[1]));
    AND3 AND2_9_inst (.A(necount[6]), .B(necount[7]), .C(necount[8]), 
        .Y(inc_10_net));
    AND3 AND2_6_inst (.A(necount[3]), .B(necount[4]), .C(necount[5]), 
        .Y(inc_5_net));
    AND2 AND2_4_inst (.A(inc_2_net), .B(necount[3]), .Y(Rcout_4_net));
    AND3 AND2_3_inst (.A(necount[0]), .B(necount[1]), .C(necount[2]), 
        .Y(inc_2_net));
    XOR2 XOR2_6_inst (.A(Rcout_8_net), .B(necount[8]), .Y(necount1[8]));
    XOR2 XOR2_1_5_inst (.A(Rcout_7_net), .B(necount[7]), .Y(
        necount1[7]));
    GND GND_i_0 (.Y(GND_0));
    AND3 AND2_11_inst (.A(inc_14_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_11_net));
    AND2 AND2_8_inst (.A(necount[6]), .B(necount[7]), .Y(inc_8_net));
    AND3 AND2_1_8_inst (.A(inc_2_net), .B(inc_5_net), .C(inc_8_net), 
        .Y(Rcout_8_net));
    XOR2 XOR2_3_inst (.A(Rcout_4_net), .B(necount[4]), .Y(necount1[4]));
    XOR2 XOR2_5_inst (.A(Rcout_6_net), .B(necount[6]), .Y(necount1[6]));
    VCC VCC_i (.Y(VCC));
    XOR2 XOR2_2_1_inst (.A(inc_1_net), .B(necount[2]), .Y(necount1[2]));
    GND GND_i (.Y(GND));
    AND3 AND2_10_inst (.A(incb_2_net), .B(necount[9]), .C(necount[10]), 
        .Y(inc_14_net));
    AND3 AND2_1_7_inst (.A(inc_2_net), .B(inc_5_net), .C(necount[6]), 
        .Y(Rcout_7_net));
    AND3 FND2_9_inst (.A(inc_12_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_10_net));
    VCC VCC_i_0 (.Y(VCC_0));
    XOR2 XOR2_7_inst (.A(Rcout_9_net), .B(necount[9]), .Y(necount1[9]));
    XOR2 XOR2_2_inst (.A(inc_2_net), .B(necount[3]), .Y(necount1[3]));
    AND2 FND2_8_inst (.A(incb_2_net), .B(necount[9]), .Y(inc_12_net));
    XOR2 FOR2_8_inst (.A(Rcout_10_net), .B(necount[10]), .Y(
        necount1[10]));
    XOR2 XOR2_9_inst (.A(Rcout_11_net), .B(necount[11]), .Y(
        necount1[11]));
    AND2 AND2_2_inst (.A(necount[0]), .B(necount[1]), .Y(inc_1_net));
    AND3 fAND2_8_inst (.A(incb_2_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_9_net));
    AND2 AND2_7_inst (.A(inc_2_net), .B(inc_5_net), .Y(Rcout_6_net));
    
endmodule


module necount_cmp_1(
       NE_NUM,
       necount,
       necount_LE_NE_1
    );
input  [11:0] NE_NUM;
input  [11:0] necount;
output necount_LE_NE_1;

    wire AND3_3_Y, XNOR2_2_Y, XNOR2_1_Y, XNOR2_10_Y, OR2A_7_Y, 
        NAND3A_4_Y, OR2A_1_Y, NAND3A_7_Y, OR2A_2_Y, OR2A_4_Y, 
        XNOR2_6_Y, XNOR2_7_Y, AO1_0_Y, NAND3A_1_Y, NAND3A_6_Y, 
        NAND3A_0_Y, NOR3A_0_Y, NAND3A_2_Y, XNOR2_0_Y, OR2A_6_Y, 
        NOR3A_1_Y, AO1C_1_Y, OR2A_3_Y, XNOR2_9_Y, AO1_1_Y, AND3_2_Y, 
        NAND3A_5_Y, XNOR2_4_Y, NOR3A_2_Y, NAND3A_3_Y, XNOR2_8_Y, 
        AND3_1_Y, XNOR2_5_Y, XNOR2_3_Y, OR2A_0_Y, NOR3A_3_Y, AND3_0_Y, 
        AND2_0_Y, OR2A_5_Y, AO1C_0_Y, XNOR2_11_Y, AO1C_2_Y, AO1C_3_Y, 
        GND, VCC, GND_0, VCC_0;
    
    OR2A OR2A_1 (.A(NE_NUM[11]), .B(necount[11]), .Y(OR2A_1_Y));
    XNOR2 XNOR2_3 (.A(necount[8]), .B(NE_NUM[8]), .Y(XNOR2_3_Y));
    NAND3A NAND3A_2 (.A(NE_NUM[4]), .B(necount[4]), .C(OR2A_0_Y), .Y(
        NAND3A_2_Y));
    NAND3A NAND3A_6 (.A(NOR3A_1_Y), .B(OR2A_6_Y), .C(NAND3A_4_Y), .Y(
        NAND3A_6_Y));
    NOR3A NOR3A_1 (.A(OR2A_1_Y), .B(AO1C_0_Y), .C(NE_NUM[9]), .Y(
        NOR3A_1_Y));
    AND3 AND3_2 (.A(XNOR2_0_Y), .B(XNOR2_11_Y), .C(XNOR2_8_Y), .Y(
        AND3_2_Y));
    AO1C AO1C_3 (.A(necount[4]), .B(NE_NUM[4]), .C(necount[3]), .Y(
        AO1C_3_Y));
    AND2 AND2_0 (.A(XNOR2_4_Y), .B(XNOR2_6_Y), .Y(AND2_0_Y));
    NOR3A NOR3A_2 (.A(OR2A_3_Y), .B(AO1C_2_Y), .C(NE_NUM[6]), .Y(
        NOR3A_2_Y));
    VCC VCC_i (.Y(VCC));
    AO1 AO1_1 (.A(AND3_2_Y), .B(NAND3A_5_Y), .C(NAND3A_0_Y), .Y(
        AO1_1_Y));
    NAND3A NAND3A_4 (.A(NE_NUM[10]), .B(necount[10]), .C(OR2A_1_Y), .Y(
        NAND3A_4_Y));
    XNOR2 XNOR2_9 (.A(necount[6]), .B(NE_NUM[6]), .Y(XNOR2_9_Y));
    NAND3A NAND3A_1 (.A(NOR3A_2_Y), .B(OR2A_4_Y), .C(NAND3A_3_Y), .Y(
        NAND3A_1_Y));
    AND3 AND3_0 (.A(XNOR2_7_Y), .B(AND3_1_Y), .C(AND2_0_Y), .Y(
        AND3_0_Y));
    OR2A OR2A_3 (.A(NE_NUM[8]), .B(necount[8]), .Y(OR2A_3_Y));
    XNOR2 XNOR2_4 (.A(necount[10]), .B(NE_NUM[10]), .Y(XNOR2_4_Y));
    OR2A OR2A_6 (.A(necount[11]), .B(NE_NUM[11]), .Y(OR2A_6_Y));
    AO1C AO1C_0 (.A(necount[10]), .B(NE_NUM[10]), .C(necount[9]), .Y(
        AO1C_0_Y));
    XNOR2 XNOR2_1 (.A(NE_NUM[10]), .B(necount[10]), .Y(XNOR2_1_Y));
    XNOR2 XNOR2_8 (.A(NE_NUM[5]), .B(necount[5]), .Y(XNOR2_8_Y));
    XNOR2 XNOR2_5 (.A(necount[7]), .B(NE_NUM[7]), .Y(XNOR2_5_Y));
    OR2A OR2A_7 (.A(necount[5]), .B(NE_NUM[5]), .Y(OR2A_7_Y));
    XNOR2 XNOR2_6 (.A(necount[11]), .B(NE_NUM[11]), .Y(XNOR2_6_Y));
    GND GND_i (.Y(GND));
    XNOR2 XNOR2_10 (.A(NE_NUM[11]), .B(necount[11]), .Y(XNOR2_10_Y));
    NOR3A NOR3A_0 (.A(OR2A_0_Y), .B(AO1C_3_Y), .C(NE_NUM[3]), .Y(
        NOR3A_0_Y));
    NAND3A NAND3A_3 (.A(NE_NUM[7]), .B(necount[7]), .C(OR2A_3_Y), .Y(
        NAND3A_3_Y));
    XNOR2 XNOR2_2 (.A(NE_NUM[9]), .B(necount[9]), .Y(XNOR2_2_Y));
    NAND3A NAND3A_5 (.A(NOR3A_3_Y), .B(OR2A_5_Y), .C(NAND3A_7_Y), .Y(
        NAND3A_5_Y));
    AND3 AND3_3 (.A(XNOR2_2_Y), .B(XNOR2_1_Y), .C(XNOR2_10_Y), .Y(
        AND3_3_Y));
    AND3 AND3_1 (.A(XNOR2_9_Y), .B(XNOR2_5_Y), .C(XNOR2_3_Y), .Y(
        AND3_1_Y));
    NAND3A NAND3A_7 (.A(NE_NUM[1]), .B(necount[1]), .C(OR2A_2_Y), .Y(
        NAND3A_7_Y));
    OR2A OR2A_4 (.A(necount[8]), .B(NE_NUM[8]), .Y(OR2A_4_Y));
    OR2A OR2A_0 (.A(NE_NUM[5]), .B(necount[5]), .Y(OR2A_0_Y));
    AO1C AO1C_1 (.A(necount[1]), .B(NE_NUM[1]), .C(necount[0]), .Y(
        AO1C_1_Y));
    XNOR2 XNOR2_11 (.A(NE_NUM[4]), .B(necount[4]), .Y(XNOR2_11_Y));
    XNOR2 XNOR2_0 (.A(NE_NUM[3]), .B(necount[3]), .Y(XNOR2_0_Y));
    OR2A OR2A_2 (.A(NE_NUM[2]), .B(necount[2]), .Y(OR2A_2_Y));
    AO1C AO1C_2 (.A(necount[7]), .B(NE_NUM[7]), .C(necount[6]), .Y(
        AO1C_2_Y));
    OR2A OR2A_5 (.A(necount[2]), .B(NE_NUM[2]), .Y(OR2A_5_Y));
    AO1 AO1_0 (.A(AND3_3_Y), .B(NAND3A_1_Y), .C(NAND3A_6_Y), .Y(
        AO1_0_Y));
    NOR3A NOR3A_3 (.A(OR2A_2_Y), .B(AO1C_1_Y), .C(NE_NUM[0]), .Y(
        NOR3A_3_Y));
    XNOR2 XNOR2_7 (.A(necount[9]), .B(NE_NUM[9]), .Y(XNOR2_7_Y));
    NAND3A NAND3A_0 (.A(NOR3A_0_Y), .B(OR2A_7_Y), .C(NAND3A_2_Y), .Y(
        NAND3A_0_Y));
    AOI1 AOI1_ALEB (.A(AND3_0_Y), .B(AO1_1_Y), .C(AO1_0_Y), .Y(
        necount_LE_NE_1));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module scalestate(
       timecount,
       scaledatain,
       strippluse,
       s_acqnum_1,
       scalechoice,
       net_45,
       timer_top_0_clk_en_scale,
       scalestate_0_dump_start,
       scalestate_0_soft_d,
       scalestate_0_rt_sw,
       net_51,
       scalestate_0_long_opentime,
       scalestate_0_s_acq,
       scalestate_0_pluse_start,
       s_acq180_c,
       scalestate_0_tetw_pluse,
       scalestate_0_dumpoff_ctr,
       top_code_0_pn_change,
       scalestate_0_dump_sustain_ctrl,
       scalestate_0_dds_conf,
       calcuinter_c,
       scalestate_0_off_test,
       scalestate_0_load_out,
       scalestate_0_pn_out,
       scalestate_0_sw_acq1,
       scalestate_0_sw_acq2,
       top_code_0_scaleload,
       timer_top_0_clk_en_scale_0,
       top_code_0_scale_rst,
       GLA
    );
output [21:0] timecount;
input  [15:0] scaledatain;
output [11:0] strippluse;
output [11:0] s_acqnum_1;
input  [4:0] scalechoice;
output net_45;
input  timer_top_0_clk_en_scale;
output scalestate_0_dump_start;
output scalestate_0_soft_d;
output scalestate_0_rt_sw;
output net_51;
output scalestate_0_long_opentime;
output scalestate_0_s_acq;
output scalestate_0_pluse_start;
output s_acq180_c;
output scalestate_0_tetw_pluse;
output scalestate_0_dumpoff_ctr;
input  top_code_0_pn_change;
output scalestate_0_dump_sustain_ctrl;
output scalestate_0_dds_conf;
output calcuinter_c;
output scalestate_0_off_test;
output scalestate_0_load_out;
output scalestate_0_pn_out;
output scalestate_0_sw_acq1;
output scalestate_0_sw_acq2;
input  top_code_0_scaleload;
input  timer_top_0_clk_en_scale_0;
input  top_code_0_scale_rst;
input  GLA;

    wire \CS_0[11]_net_1 , \CS_RNICUBC[10]_net_1 , \NS_0[8] , 
        necount_LE_NE_net_1, \CS[17]_net_1 , \CS[7]_net_1 , 
        un1_CS6_39_i_a2_2, un1_CS6_39_i_a2_1, un1_CS6_39_i_a2_0, 
        \CS[18]_net_1 , \CS_i[0]_net_1 , \timecount_18_iv_8[6] , 
        \timecount_18_iv_1[6] , \timecount_18_iv_0[6] , 
        \timecount_18_iv_6[6] , \timecount_18_iv_7[6] , 
        \CUTTIME180_TEL_m[6] , \OPENTIME_m[6] , \timecount_18_iv_4[6] , 
        \CUTTIME180_m[6] , \CUTTIME90_m[6] , \S_DUMPTIME_m[6] , 
        timecount_15_sqmuxa, \CUTTIME180_Tini[6]_net_1 , 
        \OPENTIME_TEL_m[6] , \PLUSETIME180[6]_net_1 , N_1156_i_0, 
        \PLUSETIME90_m[6] , N_1185_i_0, \DUMPTIME[6]_net_1 , 
        \ACQTIME_m[6] , \timecount_18_iv_9[7] , \timecount_18_iv_6[7] , 
        \timecount_18_iv_5[7] , \timecount_18_iv_7[7] , 
        \OPENTIME_TEL_m[7] , \CUTTIME180_Tini_m[7] , 
        \timecount_18_iv_3[7] , \S_DUMPTIME[7]_net_1 , N_1188_i_0, 
        \timecount_18_iv_2[7] , \DUMPTIME_m[7] , \ACQTIME_m[7] , 
        \timecount_18_iv_1[7] , timecount_12_sqmuxa, 
        \OPENTIME[7]_net_1 , \CUTTIME180_TEL_m[7] , N_1162_i_0, 
        \CUTTIME90[7]_net_1 , \CUTTIME180_m[7] , 
        \PLUSETIME180[7]_net_1 , \PLUSETIME90_m[7] , 
        \timecount_18_iv_8[2] , \timecount_18_iv_2[2] , 
        \S_DUMPTIME_m[2] , \timecount_18_iv_5[2] , 
        \timecount_18_iv_7[2] , \OPENTIME_TEL_m[2] , 
        \CUTTIME180_Tini_m[2] , \timecount_18_iv_3[2] , 
        \DUMPTIME_m[2] , \ACQTIME_m[2] , \timecount_18_iv_1[2] , 
        \OPENTIME[2]_net_1 , \CUTTIME180_TEL_m[2] , 
        \CUTTIME90[2]_net_1 , \CUTTIME180_m[2] , 
        \PLUSETIME180[2]_net_1 , \PLUSETIME90_m[2] , 
        timecount_18_iv_9_m1_e_9, timecount_18_iv_9_m1_e_6, 
        timecount_18_iv_9_m1_e_5, timecount_18_iv_9_m1_e_7, 
        \OPENTIME_TEL_m[9] , \CUTTIME180_Tini_m[9] , 
        timecount_18_iv_9_m1_e_3, \S_DUMPTIME[9]_net_1 , 
        timecount_18_iv_9_m1_e_2, \DUMPTIME_m[9] , \ACQTIME_m[9] , 
        timecount_18_iv_9_m1_e_1, \OPENTIME[9]_net_1 , 
        \CUTTIME180_TEL_m[9] , \CUTTIME90[9]_net_1 , \CUTTIME180_m[9] , 
        \PLUSETIME180[9]_net_1 , \PLUSETIME90_m[9] , 
        timecount_18_iv_3_m1_e_8, timecount_18_iv_3_m1_e_2, 
        \S_DUMPTIME_m[3] , timecount_18_iv_3_m1_e_5, 
        timecount_18_iv_3_m1_e_7, \OPENTIME_TEL_m[3] , 
        \CUTTIME180_Tini_m[3] , timecount_18_iv_3_m1_e_3, 
        \DUMPTIME_m[3] , \ACQTIME_m[3] , timecount_18_iv_3_m1_e_1, 
        \OPENTIME[3]_net_1 , \CUTTIME180_TEL_m[3] , 
        \CUTTIME90[3]_net_1 , \CUTTIME180_m[3] , 
        \PLUSETIME180[3]_net_1 , \PLUSETIME90_m[3] , 
        \timecount_18_iv_8[5] , \timecount_18_iv_2[5] , 
        \S_DUMPTIME_m[5] , \timecount_18_iv_5[5] , 
        \timecount_18_iv_7[5] , \OPENTIME_TEL_m[5] , 
        \CUTTIME180_Tini_m[5] , \timecount_18_iv_3[5] , 
        \DUMPTIME_m[5] , \ACQTIME_m[5] , \timecount_18_iv_1[5] , 
        \OPENTIME[5]_net_1 , \CUTTIME180_TEL_m[5] , 
        \CUTTIME90[5]_net_1 , \CUTTIME180_m[5] , 
        \PLUSETIME180[5]_net_1 , \PLUSETIME90_m[5] , 
        \timecount_18_iv_9[4] , \timecount_18_iv_6[4] , 
        \timecount_18_iv_5[4] , \timecount_18_iv_7[4] , 
        \OPENTIME_TEL_m[4] , \CUTTIME180_Tini_m[4] , 
        \timecount_18_iv_3[4] , \S_DUMPTIME[4]_net_1 , 
        \timecount_18_iv_2[4] , \DUMPTIME_m[4] , \ACQTIME_m[4] , 
        \timecount_18_iv_1[4] , \OPENTIME[4]_net_1 , 
        \CUTTIME180_TEL_m[4] , \CUTTIME90[4]_net_1 , \CUTTIME180_m[4] , 
        \PLUSETIME180[4]_net_1 , \PLUSETIME90_m[4] , 
        timecount_9_sqmuxa_m_0, \CS[13]_net_1 , 
        timecount_18_ivtt_9_m1_e_0, N_1342, \timecount_18_iv_10_8[1] , 
        \timecount_18_iv_10_1[1] , \timecount_18_iv_10_0[1] , 
        \timecount_18_iv_10_6[1] , \timecount_18_iv_10_7[1] , 
        \OPENTIME_TEL_m[1] , \CUTTIME180_Tini_m[1] , 
        \timecount_18_iv_10_3[1] , \S_DUMPTIME[1]_net_1 , 
        \timecount_18_iv_10_2[1] , \OPENTIME[1]_net_1 , 
        \CUTTIME180_TEL_m[1] , \CUTTIME90[1]_net_1 , \CUTTIME180_m[1] , 
        \PLUSETIME180[1]_net_1 , \PLUSETIME90_m[1] , 
        \DUMPTIME[1]_net_1 , \ACQTIME_m[1] , \timecount_18_iv_8[13] , 
        \timecount_18_iv_2[13] , \S_DUMPTIME_m[13] , 
        \timecount_18_iv_5[13] , \DUMPTIME_m[13] , \ACQTIME_m[13] , 
        \timecount_18_iv_1[13] , \timecount_18_iv_4[13] , 
        \CUTTIME180_Tini[13]_net_1 , \OPENTIME_TEL_m[13] , 
        \timecount_18_iv_3[13] , \OPENTIME[13]_net_1 , 
        \CUTTIME180_TEL_m[13] , \CUTTIME90[13]_net_1 , 
        \CUTTIME180_m[13] , \PLUSETIME180[13]_net_1 , 
        \PLUSETIME90_m[13] , \timecount_18_iv_8[15] , 
        \timecount_18_iv_1[15] , \timecount_18_iv_0[15] , 
        \timecount_18_iv_6[15] , \CUTTIME180_m[15] , \CUTTIME90_m[15] , 
        \S_DUMPTIME_m[15] , \timecount_18_iv_4[15] , 
        \CUTTIME180_Tini[15]_net_1 , \OPENTIME_TEL_m[15] , 
        \timecount_18_iv_3[15] , \OPENTIME[15]_net_1 , 
        \CUTTIME180_TEL_m[15] , \PLUSETIME180[15]_net_1 , 
        \PLUSETIME90_m[15] , \DUMPTIME[15]_net_1 , \ACQTIME_m[15] , 
        \timecount_18_iv_8[14] , \timecount_18_iv_1[14] , 
        \timecount_18_iv_0[14] , \timecount_18_iv_6[14] , 
        \CUTTIME180_m[14] , \CUTTIME90_m[14] , \S_DUMPTIME_m[14] , 
        \timecount_18_iv_4[14] , \CUTTIME180_Tini[14]_net_1 , 
        \OPENTIME_TEL_m[14] , \timecount_18_iv_3[14] , 
        \OPENTIME[14]_net_1 , \CUTTIME180_TEL_m[14] , 
        \PLUSETIME180[14]_net_1 , \PLUSETIME90_m[14] , 
        \DUMPTIME[14]_net_1 , \ACQTIME_m[14] , \timecount_18_iv_7[10] , 
        \OPENTIME_TEL_m[10] , \CUTTIME180_Tini_m[10] , 
        \timecount_18_iv_3[10] , \timecount_18_iv_6[10] , 
        \S_DUMPTIME[10]_net_1 , \timecount_18_iv_2[10] , 
        \timecount_18_iv_5[10] , \DUMPTIME_m[10] , \ACQTIME_m[10] , 
        \timecount_18_iv_1[10] , \OPENTIME[10]_net_1 , 
        \CUTTIME180_TEL_m[10] , \CUTTIME90[10]_net_1 , 
        \CUTTIME180_m[10] , \PLUSETIME180[10]_net_1 , 
        \PLUSETIME90_m[10] , \timecount_18_iv_8[11] , 
        \timecount_18_iv_1[11] , \timecount_18_iv_0[11] , 
        \timecount_18_iv_6[11] , \CUTTIME180_m[11] , \CUTTIME90_m[11] , 
        \S_DUMPTIME_m[11] , \timecount_18_iv_4[11] , 
        \CUTTIME180_Tini[11]_net_1 , \OPENTIME_TEL_m[11] , 
        \timecount_18_iv_3[11] , \OPENTIME[11]_net_1 , 
        \CUTTIME180_TEL_m[11] , \PLUSETIME180[11]_net_1 , 
        \PLUSETIME90_m[11] , \DUMPTIME[11]_net_1 , \ACQTIME_m[11] , 
        \timecount_18_iv_7[12] , \OPENTIME_TEL_m[12] , 
        \CUTTIME180_Tini_m[12] , \timecount_18_iv_3[12] , 
        \timecount_18_iv_6[12] , \S_DUMPTIME[12]_net_1 , 
        \timecount_18_iv_2[12] , \timecount_18_iv_5[12] , 
        \DUMPTIME_m[12] , \ACQTIME_m[12] , \timecount_18_iv_1[12] , 
        \OPENTIME[12]_net_1 , \CUTTIME180_TEL_m[12] , 
        \CUTTIME90[12]_net_1 , \CUTTIME180_m[12] , 
        \PLUSETIME180[12]_net_1 , \PLUSETIME90_m[12] , 
        \timecount_18_iv_8[8] , \timecount_18_iv_2[8] , 
        \S_DUMPTIME_m[8] , \timecount_18_iv_5[8] , \DUMPTIME_m[8] , 
        \ACQTIME_m[8] , \timecount_18_iv_1[8] , \timecount_18_iv_4[8] , 
        \CUTTIME180_Tini[8]_net_1 , \OPENTIME_TEL_m[8] , 
        \timecount_18_iv_3[8] , \OPENTIME[8]_net_1 , 
        \CUTTIME180_TEL_m[8] , \CUTTIME90[8]_net_1 , \CUTTIME180_m[8] , 
        \PLUSETIME180[8]_net_1 , \PLUSETIME90_m[8] , 
        \timecount_18_iv_7[0] , \OPENTIME_TEL_m[0] , 
        \CUTTIME180_Tini_m[0] , \timecount_18_iv_3[0] , 
        \timecount_18_iv_6[0] , \S_DUMPTIME[0]_net_1 , 
        \timecount_18_iv_2[0] , \timecount_18_iv_5[0] , 
        \DUMPTIME_m[0] , \ACQTIME_m[0] , \timecount_18_iv_1[0] , 
        timecount_14_sqmuxa, \CUTTIME180_TEL[0]_net_1 , 
        \OPENTIME_m[0] , \CUTTIME90[0]_net_1 , \CUTTIME180_m[0] , 
        \PLUSETIME180[0]_net_1 , \PLUSETIME90_m[0] , 
        \timecount_18_0_iv_2[19] , \CUTTIME180_Tini[19]_net_1 , 
        \OPENTIME_TEL_m[19] , \timecount_18_0_iv_1[19] , 
        \OPENTIME[19]_net_1 , \CUTTIME180_TEL_m[19] , 
        \timecount_18_0_iv_0[19] , \CUTTIME90[19]_net_1 , 
        \CUTTIME180_m[19] , \timecount_18_0_iv_2[17] , 
        \CUTTIME180_Tini[17]_net_1 , \OPENTIME_TEL_m[17] , 
        \timecount_18_0_iv_1[17] , \OPENTIME[17]_net_1 , 
        \CUTTIME180_TEL_m[17] , \timecount_18_0_iv_0[17] , 
        \CUTTIME90[17]_net_1 , \CUTTIME180_m[17] , 
        \timecount_18_0_iv_2[18] , \CUTTIME180_Tini[18]_net_1 , 
        \OPENTIME_TEL_m[18] , \timecount_18_0_iv_1[18] , 
        \OPENTIME[18]_net_1 , \CUTTIME180_TEL_m[18] , 
        \timecount_18_0_iv_0[18] , \CUTTIME90[18]_net_1 , 
        \CUTTIME180_m[18] , \timecount_18_0_iv_2[16] , 
        \CUTTIME180_Tini[16]_net_1 , \OPENTIME_TEL_m[16] , 
        \timecount_18_0_iv_1[16] , \OPENTIME[16]_net_1 , 
        \CUTTIME180_TEL_m[16] , \timecount_18_0_iv_0[16] , 
        \CUTTIME90[16]_net_1 , \CUTTIME180_m[16] , 
        \timecount_18_0_iv_0[20] , \CUTTIME90[20]_net_1 , 
        \CUTTIME180_TEL_m[20] , \timecount_18_0_iv_0[21] , 
        \CUTTIME90[21]_net_1 , \CUTTIME180_TEL_m[21] , 
        ACQTIME_1_sqmuxa_0_a2_0_net_1, NE_NUM_1_sqmuxa_0_a2_0_net_1, 
        un1_CS6_0, \CS[10]_net_1 , fst_lst_pulse_net_1, \CS[9]_net_1 , 
        timecount_15_sqmuxa_1, M_pulse_net_1, \CS[15]_net_1 , 
        necount_LE_M_net_1, timecount_16_sqmuxa_1, \CS_srsts_i_0[8] , 
        \CS[8]_net_1 , un1_CS_34_i_a3_0, N_1346, N_1349, 
        fst_lst_pulse8_NE_8, fst_lst_pulse8_9_i, fst_lst_pulse8_7_i, 
        fst_lst_pulse8_NE_5, fst_lst_pulse8_NE_7, fst_lst_pulse8_6_i, 
        fst_lst_pulse8_5_i, fst_lst_pulse8_NE_3, fst_lst_pulse8_NE_6, 
        fst_lst_pulse8_2_i, fst_lst_pulse8_0_i, fst_lst_pulse8_NE_1, 
        \NE_NUM[11]_net_1 , \necount[11]_net_1 , fst_lst_pulse8_10_i, 
        \NE_NUM[8]_net_1 , \necount[8]_net_1 , fst_lst_pulse8_4_i, 
        \NE_NUM[1]_net_1 , \necount[1]_net_1 , fst_lst_pulse8_3_i, 
        M_pulse8_NE_8, M_pulse8_9_i, M_pulse8_7_i, M_pulse8_NE_5, 
        M_pulse8_NE_7, M_pulse8_6_i, M_pulse8_5_i, M_pulse8_NE_3, 
        M_pulse8_NE_6, M_pulse8_2_i, M_pulse8_0_i, M_pulse8_NE_1, 
        \M_NUM[11]_net_1 , M_pulse8_10_i, \M_NUM[8]_net_1 , 
        M_pulse8_4_i, \M_NUM[1]_net_1 , M_pulse8_3_i, 
        un1_CS6_39_i_a3_1, \CS[6]_net_1 , N_1348, 
        timecount_18_iv_1_m3_e_1_1, \CS[20]_net_1 , \CS[14]_net_1 , 
        un1_CS_32_0_a3_0, un1_CS6_17_i_a3_0, \CS[4]_net_1 , 
        timecount_18_iv_9_N_2_i_0, \CS_RNITMND1[6]_net_1 , 
        timecount_18_iv_3_N_2_i_0, \timecount_RNO_2[3]_net_1 , 
        un1_timecount_5_sqmuxatt_N_6, un1_timecount_5_sqmuxa_3, 
        un1_timecount_5_sqmuxa_5, \timecount_18[1] , 
        \timecount_RNO_0[1]_net_1 , \timecount_RNO_3[1]_net_1 , 
        N_1160_i_0, \timecount_18[2] , \timecount_cnst_m[2] , 
        \timecount_18[4] , \timecount_RNO_1[4]_net_1 , 
        \timecount_18[5] , \timecount_RNO_2[5]_net_1 , 
        \timecount_18[7] , \timecount_18[16] , \timecount_18[0] , 
        \timecount_18[8] , \timecount_18[12] , \timecount_18[11] , 
        \timecount_18[10] , \timecount_18[18] , \timecount_18[14] , 
        \timecount_18[21] , \OPENTIME_TEL_m[21] , 
        \CUTTIME180_Tini_m[21] , \timecount_cnst_m[6] , N_1347, 
        \timecount_18[6] , \timecount_18[20] , \OPENTIME_TEL_m[20] , 
        \CUTTIME180_Tini_m[20] , N_1341, N_1343, N_1179, \CS[1]_net_1 , 
        un1_CS6_28, s_acqnum_1_sqmuxa, N_1278, N_1322, N_1350, 
        \CS[16]_net_1 , un1_CS6_10, intertodsp_1_sqmuxa, un1_CS6_34, 
        N_1395, sw_acq1_1_sqmuxa, N_1328, M_pulse8_NE_i_0, 
        fst_lst_pulse8_NE_i_0, un1_CS6, N_1319, \CS_RNO_1[8] , N_1323, 
        \CS[12]_net_1 , timecount_16_sqmuxa, N_1392_i, 
        \timecount_18[15] , \timecount_18[17] , NE_NUM_1_sqmuxa, N_57, 
        ACQTIME_1_sqmuxa, \timecount_18[19] , \timecount_18[13] , 
        timecount_18_iv_1_m3_e_1, un1_PLUSETIME9030_3_i_a2_0_net_1, 
        timecount_11_sqmuxa_0, N_344, N_345, N_372, un1_NS_2, N_1247, 
        N_501, N_1393, N_1253, N_507, N_1344, N_1257, N_508, N_509, 
        N_1265, N_523, N_1255, N_526, N_1243, N_527, N_511, N_1249, 
        \necount[0]_net_1 , N_512, \necount1[1] , N_515, \necount1[4] , 
        \necount[4]_net_1 , N_516, \necount1[5] , \necount[5]_net_1 , 
        N_517, \necount1[6] , \necount[6]_net_1 , N_518, \necount1[7] , 
        \necount[7]_net_1 , N_522, \necount1[11] , N_348, 
        \s_acqnum_7[0] , N_349, \s_acqnum_7[1] , N_350, 
        \s_acqnum_7[2] , N_351, \s_acqnum_7[3] , N_352, 
        \s_acqnum_7[4] , N_353, \s_acqnum_7[5] , N_354, 
        \s_acqnum_7[6] , N_355, \s_acqnum_7[7] , N_356, 
        \s_acqnum_7[8] , N_357, \s_acqnum_7[9] , N_358, 
        \s_acqnum_7[10] , N_359, \s_acqnum_7[11] , N_360, 
        \strippluse_6[0] , N_361, \strippluse_6[1] , N_362, 
        \strippluse_6[2] , N_363, \strippluse_6[3] , N_364, 
        \strippluse_6[4] , N_365, \strippluse_6[5] , N_366, 
        \strippluse_6[6] , N_367, \strippluse_6[7] , N_368, 
        \strippluse_6[8] , N_369, \strippluse_6[9] , N_370, 
        \strippluse_6[10] , N_371, \strippluse_6[11] , 
        \necount[10]_net_1 , \NE_NUM[10]_net_1 , \M_NUM[10]_net_1 , 
        \necount[9]_net_1 , \NE_NUM[9]_net_1 , \M_NUM[9]_net_1 , 
        \NE_NUM[7]_net_1 , \M_NUM[7]_net_1 , \NE_NUM[6]_net_1 , 
        \M_NUM[6]_net_1 , \NE_NUM[5]_net_1 , \M_NUM[5]_net_1 , 
        \NE_NUM[4]_net_1 , \M_NUM[4]_net_1 , \necount[3]_net_1 , 
        \NE_NUM[3]_net_1 , \M_NUM[3]_net_1 , \necount[2]_net_1 , 
        \NE_NUM[2]_net_1 , \M_NUM[2]_net_1 , \NE_NUM[0]_net_1 , 
        \M_NUM[0]_net_1 , \PLUSETIME90[2]_net_1 , \DUMPTIME[2]_net_1 , 
        \S_DUMPTIME[2]_net_1 , \OPENTIME_TEL[2]_net_1 , 
        \ACQTIME[2]_net_1 , \CUTTIME180_TEL[2]_net_1 , 
        \CUTTIME180_Tini[2]_net_1 , \CUTTIME180[2]_net_1 , 
        \PLUSETIME90[4]_net_1 , \DUMPTIME[4]_net_1 , 
        \OPENTIME_TEL[4]_net_1 , \ACQTIME[4]_net_1 , 
        \CUTTIME180_TEL[4]_net_1 , \CUTTIME180_Tini[4]_net_1 , 
        \CUTTIME180[4]_net_1 , \PLUSETIME90[5]_net_1 , 
        \DUMPTIME[5]_net_1 , \S_DUMPTIME[5]_net_1 , 
        \OPENTIME_TEL[5]_net_1 , \ACQTIME[5]_net_1 , 
        \CUTTIME180_TEL[5]_net_1 , \CUTTIME180_Tini[5]_net_1 , 
        \CUTTIME180[5]_net_1 , \OPENTIME_TEL[1]_net_1 , 
        \ACQTIME[1]_net_1 , \CUTTIME180_TEL[1]_net_1 , 
        \CUTTIME180_Tini[1]_net_1 , \CUTTIME180[1]_net_1 , 
        \DUMPTIME[7]_net_1 , \OPENTIME_TEL[7]_net_1 , 
        \ACQTIME[7]_net_1 , \CUTTIME180_TEL[7]_net_1 , 
        \CUTTIME180_Tini[7]_net_1 , \CUTTIME180[7]_net_1 , 
        \OPENTIME_TEL[8]_net_1 , \CUTTIME180[8]_net_1 , 
        \OPENTIME_TEL[16]_net_1 , \CUTTIME180_TEL[16]_net_1 , 
        \CUTTIME180[16]_net_1 , \CS_RNO[15]_net_1 , N_1309, 
        \CS_RNO[16]_net_1 , N_1310, \PLUSETIME90[0]_net_1 , 
        \DUMPTIME[0]_net_1 , \OPENTIME_TEL[0]_net_1 , 
        \OPENTIME[0]_net_1 , \ACQTIME[0]_net_1 , 
        \CUTTIME180_Tini[0]_net_1 , \CUTTIME180[0]_net_1 , 
        \DUMPTIME[3]_net_1 , \S_DUMPTIME[3]_net_1 , 
        \OPENTIME_TEL[3]_net_1 , \ACQTIME[3]_net_1 , 
        \CUTTIME180_TEL[3]_net_1 , \CUTTIME180_Tini[3]_net_1 , 
        \CUTTIME180[3]_net_1 , \DUMPTIME[8]_net_1 , 
        \S_DUMPTIME[8]_net_1 , \ACQTIME[8]_net_1 , 
        \CUTTIME180_TEL[8]_net_1 , \DUMPTIME[10]_net_1 , 
        \OPENTIME_TEL[10]_net_1 , \ACQTIME[10]_net_1 , 
        \CUTTIME180[10]_net_1 , \PLUSETIME90[11]_net_1 , 
        \S_DUMPTIME[11]_net_1 , \CUTTIME90[11]_net_1 , 
        \OPENTIME_TEL[11]_net_1 , \ACQTIME[11]_net_1 , 
        \CUTTIME180_TEL[11]_net_1 , \CUTTIME180[11]_net_1 , 
        \DUMPTIME[12]_net_1 , \OPENTIME_TEL[12]_net_1 , 
        \ACQTIME[12]_net_1 , \CUTTIME180_TEL[12]_net_1 , 
        \CUTTIME180_Tini[12]_net_1 , \CUTTIME180[12]_net_1 , 
        \S_DUMPTIME[14]_net_1 , \CUTTIME90[14]_net_1 , 
        \OPENTIME_TEL[14]_net_1 , \ACQTIME[14]_net_1 , 
        \CUTTIME180[14]_net_1 , \OPENTIME_TEL[17]_net_1 , 
        \CUTTIME180_TEL[17]_net_1 , \OPENTIME_TEL[18]_net_1 , 
        \CUTTIME180_TEL[18]_net_1 , \CUTTIME180[18]_net_1 , 
        S_DUMPTIME_1_sqmuxa, N_58, STRIPNUM180_NUM_1_sqmuxa, N_64, 
        PLUSETIME180_1_sqmuxa, N_59, PLUSETIME90_0_sqmuxa, 
        M_NUM_1_sqmuxa, DUMPTIME_1_sqmuxa, N_1320, N_246, 
        \STRIPNUM90_NUM[10]_net_1 , \STRIPNUM180_NUM[10]_net_1 , N_247, 
        \STRIPNUM90_NUM[11]_net_1 , \STRIPNUM180_NUM[11]_net_1 , N_264, 
        \ACQ90_NUM[0]_net_1 , \ACQ180_NUM[0]_net_1 , N_265, 
        \ACQ90_NUM[1]_net_1 , \ACQ180_NUM[1]_net_1 , N_266, 
        \ACQ90_NUM[2]_net_1 , \ACQ180_NUM[2]_net_1 , N_267, 
        \ACQ90_NUM[3]_net_1 , \ACQ180_NUM[3]_net_1 , N_268, 
        \ACQ90_NUM[4]_net_1 , \ACQ180_NUM[4]_net_1 , N_269, 
        \ACQ90_NUM[5]_net_1 , \ACQ180_NUM[5]_net_1 , N_270, 
        \ACQ90_NUM[6]_net_1 , \ACQ180_NUM[6]_net_1 , N_271, 
        \ACQ90_NUM[7]_net_1 , \ACQ180_NUM[7]_net_1 , N_272, 
        \ACQ90_NUM[8]_net_1 , \ACQ180_NUM[8]_net_1 , N_273, 
        \ACQ90_NUM[9]_net_1 , \ACQ180_NUM[9]_net_1 , \NS[8] , N_274, 
        \ACQ90_NUM[10]_net_1 , \ACQ180_NUM[10]_net_1 , 
        \ACQECHO_NUM[0]_net_1 , \ACQECHO_NUM[1]_net_1 , 
        \ACQECHO_NUM[2]_net_1 , \ACQECHO_NUM[3]_net_1 , 
        \ACQECHO_NUM[4]_net_1 , \ACQECHO_NUM[5]_net_1 , 
        \ACQECHO_NUM[6]_net_1 , \ACQECHO_NUM[7]_net_1 , 
        \ACQECHO_NUM[8]_net_1 , \ACQECHO_NUM[9]_net_1 , 
        \ACQECHO_NUM[10]_net_1 , N_1345, N_1351, N_244, 
        \STRIPNUM90_NUM[8]_net_1 , \STRIPNUM180_NUM[8]_net_1 , N_245, 
        \STRIPNUM90_NUM[9]_net_1 , \STRIPNUM180_NUM[9]_net_1 , N_1337, 
        \OPENTIME_TEL[21]_net_1 , \CUTTIME180_TEL[21]_net_1 , 
        \CUTTIME180_Tini[21]_net_1 , \CS[11]_net_1 , 
        \CS_RNO[14]_net_1 , N_1308, \S_DUMPTIME[6]_net_1 , 
        \CUTTIME90[6]_net_1 , \OPENTIME_TEL[6]_net_1 , 
        \OPENTIME[6]_net_1 , \ACQTIME[6]_net_1 , 
        \CUTTIME180_TEL[6]_net_1 , \CUTTIME180[6]_net_1 , un1_CS6_33, 
        N_1394, N_1276, M_pulse_RNO_net_1, dump_sustain_ctrl_RNO_net_1, 
        dds_conf_RNO_1_net_1, intertodsp_RNO_0_net_1, 
        off_test_RNO_0_net_1, dumpoff_ctr_RNO_3, load_out_RNO_net_1, 
        pn_out_RNO_net_1, \strippluse_RNO[0]_net_1 , 
        \strippluse_RNO[1]_net_1 , \strippluse_RNO[2]_net_1 , 
        \strippluse_RNO[3]_net_1 , \strippluse_RNO[4]_net_1 , 
        \strippluse_RNO[5]_net_1 , \strippluse_RNO[6]_net_1 , 
        \strippluse_RNO[7]_net_1 , \strippluse_RNO[8]_net_1 , 
        \strippluse_RNO[9]_net_1 , \strippluse_RNO[10]_net_1 , 
        \strippluse_RNO[11]_net_1 , \s_acqnum_1_RNO[0]_net_1 , 
        \s_acqnum_1_RNO[1]_net_1 , \s_acqnum_1_RNO[2]_net_1 , 
        \s_acqnum_1_RNO[3]_net_1 , \s_acqnum_1_RNO[4]_net_1 , 
        \s_acqnum_1_RNO[5]_net_1 , \s_acqnum_1_RNO[6]_net_1 , 
        \s_acqnum_1_RNO[7]_net_1 , \s_acqnum_1_RNO[8]_net_1 , 
        \s_acqnum_1_RNO[9]_net_1 , \s_acqnum_1_RNO[10]_net_1 , 
        \s_acqnum_1_RNO[11]_net_1 , \necount_RNO[1]_net_1 , 
        \necount_RNO[4]_net_1 , \necount_RNO[5]_net_1 , 
        \necount_RNO[6]_net_1 , \necount_RNO[7]_net_1 , 
        \necount_RNO[11]_net_1 , fst_lst_pulse_RNO_net_1, 
        tetw_pluse_RNO_0, sw_acq1_RNO_0_net_1, sw_acq2_RNO_3, 
        \necount_RNO[0]_net_1 , \OPENTIME_TEL[20]_net_1 , 
        \CUTTIME180_TEL[20]_net_1 , \CUTTIME180_Tini[20]_net_1 , N_236, 
        \STRIPNUM90_NUM[0]_net_1 , \STRIPNUM180_NUM[0]_net_1 , N_237, 
        \STRIPNUM90_NUM[1]_net_1 , \STRIPNUM180_NUM[1]_net_1 , N_238, 
        \STRIPNUM90_NUM[2]_net_1 , \STRIPNUM180_NUM[2]_net_1 , N_239, 
        \STRIPNUM90_NUM[3]_net_1 , \STRIPNUM180_NUM[3]_net_1 , N_240, 
        \STRIPNUM90_NUM[4]_net_1 , \STRIPNUM180_NUM[4]_net_1 , N_241, 
        \STRIPNUM90_NUM[5]_net_1 , \STRIPNUM180_NUM[5]_net_1 , N_242, 
        \STRIPNUM90_NUM[6]_net_1 , \STRIPNUM180_NUM[6]_net_1 , N_243, 
        \STRIPNUM90_NUM[7]_net_1 , \STRIPNUM180_NUM[7]_net_1 , N_275, 
        \ACQ90_NUM[11]_net_1 , \ACQ180_NUM[11]_net_1 , 
        \ACQECHO_NUM[11]_net_1 , N_1520_i, N_1552, \CS_i_RNO_1[0] , 
        N_1305, N_1263, N_1259, s_acq_RNO_0_net_1, N_505, 
        pluse_start_RNO_2, N_506, s_acq180_RNO_net_1, N_524, N_1313, 
        N_1304, \CS_RNO[20]_net_1 , \CS_RNO[10]_net_1 , soft_d_RNO_2, 
        N_346, rt_sw_RNO_4, N_347, bb_ch_RNO_net_1, N_510, 
        long_opentime_RNO_net_1, N_525, N_1296, \CS_RNO_3[1] , N_1261, 
        N_1318, N_1267, N_1340, N_504, N_1251, \CS_RNO_3[2] , N_1297, 
        \CS_RNO_3[3] , N_1298, \CS_RNO[19]_net_1 , N_1312, 
        \CS[2]_net_1 , \CS[3]_net_1 , \CS[19]_net_1 , dump_start_RNO_2, 
        \CS_RNO_1[9] , N_1303, \CS_RNO_3[5] , N_1300, \CS[5]_net_1 , 
        necount_LE_NE_RNO_net_1, necount_LE_NE_1, 
        necount_LE_M_RNO_net_1, necount_LE_M_1, N_1302, \CS_RNO_3[7] , 
        N_1301, \CS_RNO_3[6] , N_1245, \necount_RNO[10]_net_1 , N_521, 
        \necount_RNO[9]_net_1 , N_520, \necount_RNO[8]_net_1 , N_519, 
        \necount_RNO[3]_net_1 , N_514, \necount_RNO[2]_net_1 , N_513, 
        reset_out_RNO_1_net_1, N_343, \PLUSETIME90[6]_net_1 , N_1299, 
        \CS_RNO_3[4] , \PLUSETIME90[14]_net_1 , 
        \PLUSETIME90[12]_net_1 , \PLUSETIME90[10]_net_1 , 
        \CUTTIME180[9]_net_1 , \CUTTIME180_Tini[9]_net_1 , 
        \CUTTIME180_TEL[9]_net_1 , \ACQTIME[9]_net_1 , 
        \OPENTIME_TEL[9]_net_1 , \DUMPTIME[9]_net_1 , 
        \PLUSETIME90[9]_net_1 , \PLUSETIME90[8]_net_1 , 
        \PLUSETIME90[3]_net_1 , N_1307, N_1306, \CS_RNO[13]_net_1 , 
        \CS_RNO[12]_net_1 , \PLUSETIME90[7]_net_1 , 
        \PLUSETIME90[1]_net_1 , \necount1[10] , \necount1[9] , 
        \necount1[8] , \necount1[3] , \necount1[2] , N_1311, N_1289, 
        \CS_RNO[18]_net_1 , \CS_RNO[17]_net_1 , \CUTTIME180[15]_net_1 , 
        \CUTTIME180_TEL[15]_net_1 , \ACQTIME[15]_net_1 , 
        \OPENTIME_TEL[15]_net_1 , \CUTTIME90[15]_net_1 , 
        \S_DUMPTIME[15]_net_1 , \PLUSETIME90[15]_net_1 , 
        \CUTTIME180[17]_net_1 , \CUTTIME180_TEL[14]_net_1 , 
        \CUTTIME180_Tini[10]_net_1 , \CUTTIME180_TEL[10]_net_1 , 
        STRIPNUM90_NUM_1_sqmuxa, ACQ180_NUM_1_sqmuxa_1, 
        ACQECHO_NUM_1_sqmuxa, ACQ90_NUM_1_sqmuxa_1, 
        ACQ180_NUM_1_sqmuxa, N_63, ACQ90_NUM_1_sqmuxa, N_1640, N_62, 
        N_1608_i, N_1596, N_1564_i, N_1508, N_1476_i, N_1468, N_1436_i, 
        N_1428, N_1396_i, \CUTTIME180[19]_net_1 , 
        \CUTTIME180_TEL[19]_net_1 , \OPENTIME_TEL[19]_net_1 , 
        \CUTTIME180[13]_net_1 , \CUTTIME180_TEL[13]_net_1 , 
        \ACQTIME[13]_net_1 , \OPENTIME_TEL[13]_net_1 , 
        \S_DUMPTIME[13]_net_1 , \DUMPTIME[13]_net_1 , 
        \PLUSETIME90[13]_net_1 , GND, VCC, GND_0, VCC_0;
    
    DFN1E1 \DUMPTIME[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[1]_net_1 ));
    OR2B \timecount_RNO_6[8]  (.A(\S_DUMPTIME[8]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[8] ));
    DFN1E0 \CUTTIME90[2]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[2]_net_1 ));
    DFN1E1 \PLUSETIME90[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[8]_net_1 ));
    NOR3C \timecount_RNO_1[0]  (.A(\DUMPTIME_m[0] ), .B(\ACQTIME_m[0] )
        , .C(\timecount_18_iv_1[0] ), .Y(\timecount_18_iv_5[0] ));
    MX2 \s_acqnum_1_RNO_1[8]  (.A(N_272), .B(\ACQECHO_NUM[8]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[8] ));
    DFN1E1 \STRIPNUM90_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[3]_net_1 ));
    NOR2B \necount_RNO[11]  (.A(top_code_0_scale_rst), .B(N_522), .Y(
        \necount_RNO[11]_net_1 ));
    NOR2B \necount_RNO[6]  (.A(top_code_0_scale_rst), .B(N_517), .Y(
        \necount_RNO[6]_net_1 ));
    NOR2B \s_acqnum_1_RNO[7]  (.A(top_code_0_scale_rst), .B(N_355), .Y(
        \s_acqnum_1_RNO[7]_net_1 ));
    DFN1E1 \M_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[10]_net_1 ));
    OR2B \timecount_RNO_3[20]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[20]_net_1 ), .Y(\CUTTIME180_TEL_m[20] ));
    AOI1B \timecount_RNO_11[8]  (.A(\PLUSETIME180[8]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[8] ), .Y(\timecount_18_iv_1[8] )
        );
    DFN1E0 \CUTTIME180_Tini[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[4]_net_1 ));
    DFN1 \CS[11]  (.D(\CS_RNICUBC[10]_net_1 ), .CLK(GLA), .Q(
        \CS[11]_net_1 ));
    NOR3C \timecount_RNO_7[8]  (.A(\DUMPTIME_m[8] ), .B(\ACQTIME_m[8] )
        , .C(\timecount_18_iv_1[8] ), .Y(\timecount_18_iv_5[8] ));
    OR2B \timecount_RNO_4[18]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[18]_net_1 ), .Y(\CUTTIME180_m[18] ));
    OR3 \CS_RNID1N[20]  (.A(\CS[20]_net_1 ), .B(\CS[14]_net_1 ), .C(
        \CS[15]_net_1 ), .Y(timecount_18_iv_1_m3_e_1_1));
    DFN1E1 \ACQTIME[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[8]_net_1 ));
    OR2B \timecount_RNO_11[5]  (.A(N_1185_i_0), .B(\DUMPTIME[5]_net_1 )
        , .Y(\DUMPTIME_m[5] ));
    XA1A fst_lst_pulse_RNO_13 (.A(\NE_NUM[11]_net_1 ), .B(
        \necount[11]_net_1 ), .C(fst_lst_pulse8_10_i), .Y(
        fst_lst_pulse8_NE_5));
    NOR3C \timecount_RNO_1[7]  (.A(\timecount_18_iv_6[7] ), .B(
        \timecount_18_iv_5[7] ), .C(\timecount_18_iv_7[7] ), .Y(
        \timecount_18_iv_9[7] ));
    NOR2B \strippluse_RNO[6]  (.A(top_code_0_scale_rst), .B(N_366), .Y(
        \strippluse_RNO[6]_net_1 ));
    AOI1B \timecount_RNO_6[14]  (.A(N_1185_i_0), .B(
        \DUMPTIME[14]_net_1 ), .C(\ACQTIME_m[14] ), .Y(
        \timecount_18_iv_0[14] ));
    OR3C CUTTIME180_Tini_281_e (.A(N_62), .B(
        un1_PLUSETIME9030_3_i_a2_0_net_1), .C(scalechoice[0]), .Y(
        N_1596));
    NOR3C \timecount_RNO_1[6]  (.A(\CUTTIME180_TEL_m[6] ), .B(
        \OPENTIME_m[6] ), .C(\timecount_18_iv_4[6] ), .Y(
        \timecount_18_iv_7[6] ));
    DFN1E1 \timecount[14]  (.D(\timecount_18[14] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[14]));
    DFN1E0 \CUTTIME180_TEL[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[8]_net_1 ));
    NOR3B un1_PLUSETIME9030_4_i_a2_0 (.A(top_code_0_scaleload), .B(
        scalechoice[1]), .C(scalechoice[4]), .Y(N_57));
    OR2B \timecount_RNO_1[20]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[20]_net_1 ), .Y(\CUTTIME180_Tini_m[20] ));
    DFN1 \strippluse[10]  (.D(\strippluse_RNO[10]_net_1 ), .CLK(GLA), 
        .Q(strippluse[10]));
    OR3C \timecount_RNO_0[20]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[20]_net_1 ), .Y(
        \OPENTIME_TEL_m[20] ));
    OR3C \timecount_RNO_5[17]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[17]_net_1 ), .Y(
        \OPENTIME_TEL_m[17] ));
    AOI1B \timecount_RNO_2[21]  (.A(N_1162_i_0), .B(
        \CUTTIME90[21]_net_1 ), .C(\CUTTIME180_TEL_m[21] ), .Y(
        \timecount_18_0_iv_0[21] ));
    MX2 \s_acqnum_1_RNO_0[7]  (.A(\s_acqnum_7[7] ), .B(s_acqnum_1[7]), 
        .S(un1_CS6_28), .Y(N_355));
    OR2B \timecount_RNO_12[8]  (.A(\PLUSETIME90[8]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[8] ));
    OR3C \timecount_RNO[13]  (.A(\timecount_18_iv_4[13] ), .B(
        \timecount_18_iv_3[13] ), .C(\timecount_18_iv_8[13] ), .Y(
        \timecount_18[13] ));
    MX2C \CS_RNO_0[15]  (.A(\CS[15]_net_1 ), .B(\CS[14]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1309));
    OR2 \timecount_RNO_2[5]  (.A(\CS_RNITMND1[6]_net_1 ), .B(N_1337), 
        .Y(\timecount_RNO_2[5]_net_1 ));
    DFN1 \strippluse[8]  (.D(\strippluse_RNO[8]_net_1 ), .CLK(GLA), .Q(
        strippluse[8]));
    OR2B \timecount_RNO_11[1]  (.A(\PLUSETIME90[1]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[1] ));
    NOR2B pluse_start_RNO (.A(top_code_0_scale_rst), .B(N_506), .Y(
        pluse_start_RNO_2));
    DFN1E0 \CUTTIME180_TEL[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[13]_net_1 ));
    OR2B \timecount_RNO_12[15]  (.A(\S_DUMPTIME[15]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[15] ));
    OR2B \timecount_RNO_10[4]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[4]_net_1 ), .Y(\CUTTIME180_Tini_m[4] ));
    OR2 un1_PLUSETIME9030_3_i_a2_0 (.A(scalechoice[3]), .B(
        scalechoice[2]), .Y(N_58));
    DFN1E1 \timecount[12]  (.D(\timecount_18[12] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[12]));
    MX2 \s_acqnum_1_RNO_1[9]  (.A(N_273), .B(\ACQECHO_NUM[9]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[9] ));
    DFN1E0 \CUTTIME180[2]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[2]_net_1 ));
    DFN1E1 \timecount[13]  (.D(\timecount_18[13] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[13]));
    MX2 fst_lst_pulse_RNO_0 (.A(fst_lst_pulse8_NE_i_0), .B(
        fst_lst_pulse_net_1), .S(N_1255), .Y(N_523));
    DFN1E0 \CUTTIME90[20]  (.D(scaledatain[4]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[20]_net_1 ));
    OR2B bb_ch_RNO_1 (.A(timer_top_0_clk_en_scale_0), .B(N_1347), .Y(
        N_1261));
    DFN1E1 \ACQ180_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[7]_net_1 ));
    NOR2B \s_acqnum_1_RNO[5]  (.A(top_code_0_scale_rst), .B(N_353), .Y(
        \s_acqnum_1_RNO[5]_net_1 ));
    DFN1E1 \ACQECHO_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[11]_net_1 ));
    OR2B \timecount_RNO_7[3]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[3]_net_1 ), .Y(\CUTTIME180_Tini_m[3] ));
    DFN1E1 \ACQ180_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[4]_net_1 ));
    DFN1E1 \M_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[1]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[3]_net_1 ));
    OR2B \CS_RNI4897[13]  (.A(N_1278), .B(\CS[13]_net_1 ), .Y(N_1249));
    MX2 \strippluse_RNO_0[11]  (.A(\strippluse_6[11] ), .B(
        strippluse[11]), .S(un1_CS6_28), .Y(N_371));
    DFN1E0 \CUTTIME180[16]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1428), 
        .Q(\CUTTIME180[16]_net_1 ));
    OR2 \CS_RNIR8F[12]  (.A(\CS[13]_net_1 ), .B(\CS[12]_net_1 ), .Y(
        N_1348));
    DFN1 \CS[4]  (.D(\CS_RNO_3[4] ), .CLK(GLA), .Q(\CS[4]_net_1 ));
    NOR3C \timecount_RNO_0[4]  (.A(\timecount_18_iv_6[4] ), .B(
        \timecount_18_iv_5[4] ), .C(\timecount_18_iv_7[4] ), .Y(
        \timecount_18_iv_9[4] ));
    OA1C \CS_RNI1K67[18]  (.A(\CS[17]_net_1 ), .B(necount_LE_NE_net_1), 
        .C(\CS[18]_net_1 ), .Y(N_1394));
    OR3C \timecount_RNO_5[0]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[0]_net_1 ), .Y(
        \ACQTIME_m[0] ));
    DFN1E1 \NE_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[7]_net_1 ));
    OR2B \timecount_RNO_12[0]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[0]_net_1 ), .Y(\OPENTIME_m[0] ));
    DFN1E1 \timecount[19]  (.D(\timecount_18[19] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[19]));
    DFN1E0 \CUTTIME180_TEL[16]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[16]_net_1 ));
    OR3C \timecount_RNO_3[13]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[13]_net_1 ), .Y(
        \OPENTIME_TEL_m[13] ));
    DFN1E1 \timecount[6]  (.D(\timecount_18[6] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[6]));
    MX2 s_acq180_RNO_0 (.A(\CS[9]_net_1 ), .B(s_acq180_c), .S(un1_CS6), 
        .Y(N_524));
    DFN1E1 \ACQTIME[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[15]_net_1 ));
    DFN1E1 \DUMPTIME[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[8]_net_1 ));
    DFN1 dumpoff_ctr (.D(dumpoff_ctr_RNO_3), .CLK(GLA), .Q(
        scalestate_0_dumpoff_ctr));
    AOI1B \timecount_RNO_8[2]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[2]_net_1 ), .C(\CUTTIME180_TEL_m[2] ), .Y(
        \timecount_18_iv_3[2] ));
    NOR2A \CS_RNO[16]  (.A(top_code_0_scale_rst), .B(N_1310), .Y(
        \CS_RNO[16]_net_1 ));
    MX2 pn_out_RNO_0 (.A(un1_NS_2), .B(scalestate_0_pn_out), .S(N_1247)
        , .Y(N_372));
    MX2 s_acq180_RNO_2 (.A(\CS[10]_net_1 ), .B(fst_lst_pulse_net_1), 
        .S(\CS[9]_net_1 ), .Y(un1_CS6_0));
    NOR2 \strippluse_RNO_1[5]  (.A(N_241), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[5] ));
    DFN1 \strippluse[9]  (.D(\strippluse_RNO[9]_net_1 ), .CLK(GLA), .Q(
        strippluse[9]));
    OR2B \timecount_RNO_10[2]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[2]_net_1 ), .Y(\CUTTIME180_m[2] ));
    OR2B \timecount_RNO_9[6]  (.A(\PLUSETIME90[6]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[6] ));
    OR2B \timecount_RNO[4]  (.A(\timecount_18_iv_9[4] ), .B(
        \timecount_RNO_1[4]_net_1 ), .Y(\timecount_18[4] ));
    MX2 \s_acqnum_1_RNO_1[5]  (.A(N_269), .B(\ACQECHO_NUM[5]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[5] ));
    AOI1B \timecount_RNO_2[20]  (.A(N_1162_i_0), .B(
        \CUTTIME90[20]_net_1 ), .C(\CUTTIME180_TEL_m[20] ), .Y(
        \timecount_18_0_iv_0[20] ));
    DFN1 \CS_0[11]  (.D(\CS_RNICUBC[10]_net_1 ), .CLK(GLA), .Q(
        \CS_0[11]_net_1 ));
    AOI1B \timecount_RNO_5[15]  (.A(\PLUSETIME180[15]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[15] ), .Y(
        \timecount_18_iv_1[15] ));
    OR2B \timecount_RNO_10[11]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[11]_net_1 ), .Y(\CUTTIME180_m[11] ));
    NOR3B S_DUMPTIME_1_sqmuxa_0_a2 (.A(scalechoice[0]), .B(N_57), .C(
        N_58), .Y(S_DUMPTIME_1_sqmuxa));
    DFN1E1 \ACQ180_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[11]_net_1 ));
    MX2C \strippluse_RNO_2[0]  (.A(\STRIPNUM90_NUM[0]_net_1 ), .B(
        \STRIPNUM180_NUM[0]_net_1 ), .S(\NS[8] ), .Y(N_236));
    DFN1E0 \CUTTIME90[21]  (.D(scaledatain[5]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[21]_net_1 ));
    NOR2 \strippluse_RNO_1[7]  (.A(N_243), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[7] ));
    MX2C \CS_RNO_0[2]  (.A(\CS[2]_net_1 ), .B(\CS[1]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1297));
    NOR2B \strippluse_RNO[7]  (.A(top_code_0_scale_rst), .B(N_367), .Y(
        \strippluse_RNO[7]_net_1 ));
    OR2A reset_out_RNO_3 (.A(\CS_i[0]_net_1 ), .B(\CS[6]_net_1 ), .Y(
        un1_CS_32_0_a3_0));
    DFN1E0 \CUTTIME90[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[15]_net_1 ));
    MX2C \CS_RNO_0[4]  (.A(\CS[4]_net_1 ), .B(\CS[19]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1299));
    OR2B \timecount_RNO_11[11]  (.A(N_1162_i_0), .B(
        \CUTTIME90[11]_net_1 ), .Y(\CUTTIME90_m[11] ));
    OR2B \timecount_RNO_3[18]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[18]_net_1 ), .Y(\CUTTIME180_TEL_m[18] ));
    DFN1 \s_acqnum_1[11]  (.D(\s_acqnum_1_RNO[11]_net_1 ), .CLK(GLA), 
        .Q(s_acqnum_1[11]));
    AOI1B \timecount_RNO_3[2]  (.A(N_1162_i_0), .B(
        \CUTTIME90[2]_net_1 ), .C(\CUTTIME180_m[2] ), .Y(
        \timecount_18_iv_2[2] ));
    MX2A sw_acq2_RNO_0 (.A(N_1348), .B(scalestate_0_sw_acq2), .S(
        un1_CS6_34), .Y(N_344));
    DFN1E0 \OPENTIME_TEL[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[1]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[3]_net_1 ));
    AOI1B \timecount_RNO_0[16]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[16]_net_1 ), .C(\CUTTIME180_TEL_m[16] ), .Y(
        \timecount_18_0_iv_1[16] ));
    DFN1E1 \PLUSETIME90[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[6]_net_1 ));
    DFN1E0 \CUTTIME180[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[14]_net_1 ));
    NOR3C M_pulse_RNO_4 (.A(M_pulse8_9_i), .B(M_pulse8_7_i), .C(
        M_pulse8_NE_5), .Y(M_pulse8_NE_8));
    DFN1E0 \OPENTIME[13]  (.D(scaledatain[13]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[13]_net_1 ));
    OR3C \timecount_RNO[2]  (.A(\timecount_18_iv_8[2] ), .B(
        \timecount_18_iv_7[2] ), .C(\timecount_cnst_m[2] ), .Y(
        \timecount_18[2] ));
    OR2B \timecount_RNO_13[3]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[3]_net_1 ), .Y(\CUTTIME180_TEL_m[3] ));
    AO1 \timecount_RNO_1[4]  (.A(top_code_0_scale_rst), .B(N_1341), .C(
        \CS_RNITMND1[6]_net_1 ), .Y(\timecount_RNO_1[4]_net_1 ));
    MX2C \strippluse_RNO_2[11]  (.A(\STRIPNUM90_NUM[11]_net_1 ), .B(
        \STRIPNUM180_NUM[11]_net_1 ), .S(\NS_0[8] ), .Y(N_247));
    DFN1E1 \STRIPNUM90_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[0]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[10]_net_1 ));
    MX2C \CS_RNO_0[6]  (.A(\CS[6]_net_1 ), .B(\CS[5]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1301));
    NOR3A STRIPNUM180_NUM_1_sqmuxa_0_a2 (.A(N_64), .B(N_58), .C(
        scalechoice[0]), .Y(STRIPNUM180_NUM_1_sqmuxa));
    DFN1E1 \PLUSETIME180[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[0]_net_1 ));
    DFN1E1 \timecount[0]  (.D(\timecount_18[0] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[0]));
    DFN1E0 \CUTTIME180[5]  (.D(scaledatain[5]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[5]_net_1 ));
    DFN1 \s_acqnum_1[4]  (.D(\s_acqnum_1_RNO[4]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[4]));
    AOI1B \timecount_RNO_5[14]  (.A(\PLUSETIME180[14]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[14] ), .Y(
        \timecount_18_iv_1[14] ));
    DFN1E0 \CUTTIME180_TEL[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[1]_net_1 ));
    AOI1B \timecount_RNO_0[8]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[8]_net_1 ), .C(\OPENTIME_TEL_m[8] ), .Y(
        \timecount_18_iv_4[8] ));
    DFN1 sw_acq1 (.D(sw_acq1_RNO_0_net_1), .CLK(GLA), .Q(
        scalestate_0_sw_acq1));
    AOI1B \timecount_RNO_5[7]  (.A(N_1162_i_0), .B(
        \CUTTIME90[7]_net_1 ), .C(\CUTTIME180_m[7] ), .Y(
        \timecount_18_iv_2[7] ));
    AOI1B \timecount_RNO_1[19]  (.A(N_1162_i_0), .B(
        \CUTTIME90[19]_net_1 ), .C(\CUTTIME180_m[19] ), .Y(
        \timecount_18_0_iv_0[19] ));
    DFN1E1 \timecount[10]  (.D(\timecount_18[10] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[10]));
    OR2B \timecount_RNO_10[12]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[12]_net_1 ), .Y(\CUTTIME180_m[12] ));
    DFN1E1 \DUMPTIME[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[4]_net_1 ));
    NOR2B \strippluse_RNO[1]  (.A(top_code_0_scale_rst), .B(N_361), .Y(
        \strippluse_RNO[1]_net_1 ));
    DFN1E1 \DUMPTIME[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[2]_net_1 ));
    NOR2A \CS_RNO[2]  (.A(top_code_0_scale_rst), .B(N_1297), .Y(
        \CS_RNO_3[2] ));
    OR2B \timecount_RNO_14[3]  (.A(\PLUSETIME90[3]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[3] ));
    OR2B \timecount_RNO_11[12]  (.A(\PLUSETIME90[12]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[12] ));
    NOR3C \timecount_RNO_2[13]  (.A(\timecount_18_iv_2[13] ), .B(
        \S_DUMPTIME_m[13] ), .C(\timecount_18_iv_5[13] ), .Y(
        \timecount_18_iv_8[13] ));
    DFN1E0 \CUTTIME90[16]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[16]_net_1 ));
    NOR2B dump_start_RNO (.A(top_code_0_scale_rst), .B(N_504), .Y(
        dump_start_RNO_2));
    NOR2A \CS_RNO[20]  (.A(top_code_0_scale_rst), .B(N_1313), .Y(
        \CS_RNO[20]_net_1 ));
    OR2A \CS_RNIN78E[18]  (.A(N_1278), .B(N_1394), .Y(N_1276));
    NOR3C \timecount_RNO_7[13]  (.A(\DUMPTIME_m[13] ), .B(
        \ACQTIME_m[13] ), .C(\timecount_18_iv_1[13] ), .Y(
        \timecount_18_iv_5[13] ));
    NOR2 \strippluse_RNO_1[8]  (.A(N_244), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[8] ));
    MX2 \s_acqnum_1_RNO_1[11]  (.A(N_275), .B(\ACQECHO_NUM[11]_net_1 ), 
        .S(\CS[11]_net_1 ), .Y(\s_acqnum_7[11] ));
    OR3C \timecount_RNO_6[5]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[5]_net_1 ), .Y(
        \OPENTIME_TEL_m[5] ));
    DFN1E1 \ACQ180_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[1]_net_1 ));
    OA1C \CS_RNO[8]  (.A(timer_top_0_clk_en_scale_0), .B(\NS_0[8] ), 
        .C(\CS_srsts_i_0[8] ), .Y(\CS_RNO_1[8] ));
    DFN1E1 \PLUSETIME180[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[3]_net_1 ));
    DFN1E1 \M_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[3]_net_1 ));
    NOR3C \timecount_RNO_0[2]  (.A(\timecount_18_iv_2[2] ), .B(
        \S_DUMPTIME_m[2] ), .C(\timecount_18_iv_5[2] ), .Y(
        \timecount_18_iv_8[2] ));
    OR3C \timecount_RNO[0]  (.A(\timecount_18_iv_6[0] ), .B(
        \timecount_18_iv_5[0] ), .C(\timecount_18_iv_7[0] ), .Y(
        \timecount_18[0] ));
    OR3A CUTTIME180_TEL_243_e (.A(un1_PLUSETIME9030_3_i_a2_0_net_1), 
        .B(N_58), .C(scalechoice[0]), .Y(N_1520_i));
    DFN1E1 \ACQTIME[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[3]_net_1 ));
    NOR2 \strippluse_RNO_1[2]  (.A(N_238), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[2] ));
    DFN1E0 \CUTTIME90[4]  (.D(scaledatain[4]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[4]_net_1 ));
    NOR3B un1_PLUSETIME9030_1_i_a2_1 (.A(top_code_0_scaleload), .B(
        scalechoice[4]), .C(scalechoice[1]), .Y(N_64));
    DFN1E1 \STRIPNUM90_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[7]_net_1 ));
    AOI1B \timecount_RNO_2[18]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[18]_net_1 ), .C(\OPENTIME_TEL_m[18] ), .Y(
        \timecount_18_0_iv_2[18] ));
    DFN1 \s_acqnum_1[2]  (.D(\s_acqnum_1_RNO[2]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[2]));
    AO1C \timecount_RNO[9]  (.A(\CS_RNITMND1[6]_net_1 ), .B(
        timecount_18_ivtt_9_m1_e_0), .C(timecount_18_iv_9_m1_e_9), .Y(
        timecount_18_iv_9_N_2_i_0));
    DFN1E0 \OPENTIME_TEL[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[6]_net_1 ));
    DFN1E1 \timecount[16]  (.D(\timecount_18[16] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[16]));
    DFN1E0 \OPENTIME[19]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1468), 
        .Q(\OPENTIME[19]_net_1 ));
    MX2C \CS_RNI2OR7[10]  (.A(\CS[11]_net_1 ), .B(\CS[10]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1305));
    AOI1B \timecount_RNO_7[1]  (.A(\PLUSETIME180[1]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[1] ), .Y(
        \timecount_18_iv_10_1[1] ));
    NOR2B s_acq180_RNO (.A(top_code_0_scale_rst), .B(N_524), .Y(
        s_acq180_RNO_net_1));
    DFN1E0 \OPENTIME[9]  (.D(scaledatain[9]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[9]_net_1 ));
    NOR2B \strippluse_RNO[2]  (.A(top_code_0_scale_rst), .B(N_362), .Y(
        \strippluse_RNO[2]_net_1 ));
    DFN1 pluse_start (.D(pluse_start_RNO_2), .CLK(GLA), .Q(
        scalestate_0_pluse_start));
    DFN1E1 \ACQTIME[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[1]_net_1 ));
    OR2B \timecount_RNO_15[5]  (.A(\PLUSETIME90[5]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[5] ));
    OA1 \timecount_RNO_0[7]  (.A(\CS[13]_net_1 ), .B(\NS_0[8] ), .C(
        top_code_0_scale_rst), .Y(timecount_9_sqmuxa_m_0));
    DFN1E0 \OPENTIME_TEL[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[5]_net_1 ));
    DFN1E0 \OPENTIME_TEL[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[3]_net_1 ));
    DFN1E1 \PLUSETIME180[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[8]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[6]_net_1 ));
    AOI1B \timecount_RNO_13[5]  (.A(\PLUSETIME180[5]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[5] ), .Y(\timecount_18_iv_1[5] )
        );
    DFN1E1 \ACQTIME[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[6]_net_1 ));
    MX2 s_acq_RNO_0 (.A(N_1342), .B(scalestate_0_s_acq), .S(N_1259), 
        .Y(N_505));
    DFN1 fst_lst_pulse (.D(fst_lst_pulse_RNO_net_1), .CLK(GLA), .Q(
        fst_lst_pulse_net_1));
    NOR2 \CS_RNIUUGC[2]  (.A(\CS[8]_net_1 ), .B(\CS[2]_net_1 ), .Y(
        N_1345));
    NOR2 \strippluse_RNO_1[9]  (.A(N_245), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[9] ));
    DFN1 \CS[12]  (.D(\CS_RNO[12]_net_1 ), .CLK(GLA), .Q(
        \CS[12]_net_1 ));
    DFN1E1 \DUMPTIME[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[3]_net_1 ));
    OR3C \timecount_RNO_9[15]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[15]_net_1 ), .Y(
        \ACQTIME_m[15] ));
    MX2 bb_ch_RNO_0 (.A(N_1320), .B(net_51), .S(N_1261), .Y(N_510));
    MX2 \s_acqnum_1_RNO_0[1]  (.A(\s_acqnum_7[1] ), .B(s_acqnum_1[1]), 
        .S(un1_CS6_28), .Y(N_349));
    NOR3C fst_lst_pulse_RNO_1 (.A(fst_lst_pulse8_NE_7), .B(
        fst_lst_pulse8_NE_6), .C(fst_lst_pulse8_NE_8), .Y(
        fst_lst_pulse8_NE_i_0));
    OR2B \timecount_RNO_10[3]  (.A(N_1185_i_0), .B(\DUMPTIME[3]_net_1 )
        , .Y(\DUMPTIME_m[3] ));
    AO1B \CS_RNIM93J[18]  (.A(timer_top_0_clk_en_scale_0), .B(N_1394), 
        .C(top_code_0_scale_rst), .Y(un1_CS6_33));
    NOR3C \timecount_RNO_3[7]  (.A(\DUMPTIME_m[7] ), .B(\ACQTIME_m[7] )
        , .C(\timecount_18_iv_1[7] ), .Y(\timecount_18_iv_5[7] ));
    OR2B \timecount_RNO_8[11]  (.A(\PLUSETIME90[11]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[11] ));
    DFN1E0 \OPENTIME_TEL[21]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[21]_net_1 ));
    MX2 \necount_RNO_0[11]  (.A(\necount1[11] ), .B(
        \necount[11]_net_1 ), .S(N_1249), .Y(N_522));
    OR2B \timecount_RNO_12[10]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[10]_net_1 ), .Y(\CUTTIME180_TEL_m[10] ));
    OAI1 \timecount_RNO_3[1]  (.A(N_1341), .B(timecount_18_iv_1_m3_e_1)
        , .C(top_code_0_scale_rst), .Y(\timecount_RNO_3[1]_net_1 ));
    DFN1 rt_sw (.D(rt_sw_RNO_4), .CLK(GLA), .Q(scalestate_0_rt_sw));
    DFN1E1 \timecount[2]  (.D(\timecount_18[2] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[2]));
    NOR3C fst_lst_pulse_RNO_4 (.A(fst_lst_pulse8_9_i), .B(
        fst_lst_pulse8_7_i), .C(fst_lst_pulse8_NE_5), .Y(
        fst_lst_pulse8_NE_8));
    DFN1E1 \S_DUMPTIME[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[14]_net_1 ));
    NOR3B \CS_RNIDRV5[12]  (.A(\CS[12]_net_1 ), .B(
        top_code_0_scale_rst), .C(necount_LE_M_net_1), .Y(
        timecount_12_sqmuxa));
    MX2 \s_acqnum_1_RNO_2[4]  (.A(\ACQ90_NUM[4]_net_1 ), .B(
        \ACQ180_NUM[4]_net_1 ), .S(\NS_0[8] ), .Y(N_268));
    DFN1E1 \ACQ180_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[0]_net_1 ));
    OR3A OPENTIME_217_e (.A(scalechoice[0]), .B(N_63), .C(
        scalechoice[2]), .Y(N_1468));
    DFN1E1 \NE_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[3]_net_1 ));
    DFN1 \s_acqnum_1[7]  (.D(\s_acqnum_1_RNO[7]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[7]));
    NOR3C \timecount_RNO_0[6]  (.A(\timecount_18_iv_1[6] ), .B(
        \timecount_18_iv_0[6] ), .C(\timecount_18_iv_6[6] ), .Y(
        \timecount_18_iv_8[6] ));
    OR2B \timecount_RNO_14[4]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[4]_net_1 ), .Y(\CUTTIME180_TEL_m[4] ));
    AOI1B \timecount_RNO_0[11]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[11]_net_1 ), .C(\OPENTIME_TEL_m[11] ), .Y(
        \timecount_18_iv_4[11] ));
    DFN1 \s_acqnum_1[8]  (.D(\s_acqnum_1_RNO[8]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[8]));
    OAI1 dump_sustain_ctrl_RNO_1 (.A(\CS[11]_net_1 ), .B(
        \CS[13]_net_1 ), .C(N_1278), .Y(N_1243));
    DFN1E1 \STRIPNUM90_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[5]_net_1 ));
    DFN1E1 \NE_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[6]_net_1 ));
    OR2B \timecount_RNO_9[2]  (.A(N_1345), .B(N_1343), .Y(N_1328));
    OR3C \timecount_RNO_9[14]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[14]_net_1 ), .Y(
        \ACQTIME_m[14] ));
    DFN1E0 \OPENTIME_TEL[16]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[16]_net_1 ));
    NOR2A \CS_RNO[9]  (.A(top_code_0_scale_rst), .B(N_1303), .Y(
        \CS_RNO_1[9] ));
    DFN1E1 \PLUSETIME180[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[9]_net_1 ));
    DFN1 tetw_pluse (.D(tetw_pluse_RNO_0), .CLK(GLA), .Q(
        scalestate_0_tetw_pluse));
    MX2 \s_acqnum_1_RNO_2[2]  (.A(\ACQ90_NUM[2]_net_1 ), .B(
        \ACQ180_NUM[2]_net_1 ), .S(\NS_0[8] ), .Y(N_266));
    NOR2B \strippluse_RNO[11]  (.A(top_code_0_scale_rst), .B(N_371), 
        .Y(\strippluse_RNO[11]_net_1 ));
    OR2B \timecount_RNO_13[7]  (.A(\PLUSETIME90[7]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[7] ));
    OA1 \CS_RNO[18]  (.A(\CS[18]_net_1 ), .B(N_1289), .C(
        top_code_0_scale_rst), .Y(\CS_RNO[18]_net_1 ));
    NOR2 \strippluse_RNO_1[0]  (.A(N_236), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[0] ));
    DFN1E1 \PLUSETIME90[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[7]_net_1 ));
    NOR2B necount_LE_NE_RNO (.A(top_code_0_scale_rst), .B(
        necount_LE_NE_1), .Y(necount_LE_NE_RNO_net_1));
    DFN1 load_out (.D(load_out_RNO_net_1), .CLK(GLA), .Q(
        scalestate_0_load_out));
    DFN1E1 \ACQECHO_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[10]_net_1 ));
    DFN1E0 \OPENTIME[17]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1468), 
        .Q(\OPENTIME[17]_net_1 ));
    AOI1B \timecount_RNO_8[3]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[3]_net_1 ), .C(\CUTTIME180_TEL_m[3] ), .Y(
        timecount_18_iv_3_m1_e_3));
    OR2A sw_acq2_RNO (.A(top_code_0_scale_rst), .B(N_344), .Y(
        sw_acq2_RNO_3));
    DFN1E0 \OPENTIME_TEL[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[13]_net_1 ));
    OR3A \CS_RNI9VUJ[13]  (.A(N_1343), .B(\CS[13]_net_1 ), .C(
        \NS_0[8] ), .Y(N_1341));
    NOR3C \timecount_RNO_1[12]  (.A(\DUMPTIME_m[12] ), .B(
        \ACQTIME_m[12] ), .C(\timecount_18_iv_1[12] ), .Y(
        \timecount_18_iv_5[12] ));
    OR2B \timecount_RNO_4[3]  (.A(\S_DUMPTIME[3]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[3] ));
    MX2 \s_acqnum_1_RNO_2[1]  (.A(\ACQ90_NUM[1]_net_1 ), .B(
        \ACQ180_NUM[1]_net_1 ), .S(\NS_0[8] ), .Y(N_265));
    OR3C \timecount_RNO_5[16]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[16]_net_1 ), .Y(
        \OPENTIME_TEL_m[16] ));
    MX2 M_pulse_RNO_0 (.A(M_pulse8_NE_i_0), .B(M_pulse_net_1), .S(
        N_1255), .Y(N_527));
    OAI1 load_out_RNO_1 (.A(N_1351), .B(N_1393), .C(N_1278), .Y(N_1253)
        );
    NOR2 \CS_RNIPVF6[4]  (.A(\CS[10]_net_1 ), .B(\CS[4]_net_1 ), .Y(
        N_1346));
    OAI1 dds_conf_RNO_1 (.A(N_1344), .B(N_1347), .C(N_1278), .Y(N_1265)
        );
    NOR2A \CS_RNO[17]  (.A(top_code_0_scale_rst), .B(N_1311), .Y(
        \CS_RNO[17]_net_1 ));
    NOR2A NE_NUM_1_sqmuxa_0_a2_0 (.A(scalechoice[0]), .B(
        scalechoice[2]), .Y(NE_NUM_1_sqmuxa_0_a2_0_net_1));
    OR2B \timecount_RNO_8[10]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[10]_net_1 ), .Y(\CUTTIME180_Tini_m[10] ));
    DFN1E1 \DUMPTIME[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[6]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[8]_net_1 ));
    NOR3B M_NUM_1_sqmuxa_0_a2 (.A(scalechoice[0]), .B(N_64), .C(N_58), 
        .Y(M_NUM_1_sqmuxa));
    DFN1E0 \CUTTIME180[1]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[1]_net_1 ));
    AOI1B \timecount_RNO_6[11]  (.A(N_1185_i_0), .B(
        \DUMPTIME[11]_net_1 ), .C(\ACQTIME_m[11] ), .Y(
        \timecount_18_iv_0[11] ));
    MX2 \strippluse_RNO_0[6]  (.A(\strippluse_6[6] ), .B(strippluse[6])
        , .S(un1_CS6_28), .Y(N_366));
    DFN1E0 \CUTTIME180_Tini[16]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[16]_net_1 ));
    AOI1B \timecount_RNO_2[7]  (.A(\S_DUMPTIME[7]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_2[7] ), .Y(
        \timecount_18_iv_6[7] ));
    MX2 \necount_RNO_0[2]  (.A(\necount1[2] ), .B(\necount[2]_net_1 ), 
        .S(N_1249), .Y(N_513));
    OR2B \timecount_RNO_10[9]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[9]_net_1 ), .Y(\CUTTIME180_Tini_m[9] ));
    DFN1E0 \OPENTIME_TEL[17]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[17]_net_1 ));
    XNOR2 fst_lst_pulse_RNO_16 (.A(\necount[10]_net_1 ), .B(
        \NE_NUM[10]_net_1 ), .Y(fst_lst_pulse8_10_i));
    OR2B \timecount_RNO_14[7]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[7]_net_1 ), .Y(\CUTTIME180_TEL_m[7] ));
    DFN1 \CS[17]  (.D(\CS_RNO[17]_net_1 ), .CLK(GLA), .Q(
        \CS[17]_net_1 ));
    AOI1B \timecount_RNO_8[1]  (.A(N_1185_i_0), .B(\DUMPTIME[1]_net_1 )
        , .C(\ACQTIME_m[1] ), .Y(\timecount_18_iv_10_0[1] ));
    DFN1E1 \timecount[20]  (.D(\timecount_18[20] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[20]));
    OR2 \CS_RNI2DF[19]  (.A(\CS[20]_net_1 ), .B(\CS[19]_net_1 ), .Y(
        N_1344));
    OR2B \timecount_RNO_7[6]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[6]_net_1 ), .Y(\OPENTIME_m[6] ));
    XNOR2 M_pulse_RNO_14 (.A(\necount[4]_net_1 ), .B(\M_NUM[4]_net_1 ), 
        .Y(M_pulse8_4_i));
    AOI1B \timecount_RNO_0[10]  (.A(\S_DUMPTIME[10]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_2[10] ), .Y(
        \timecount_18_iv_6[10] ));
    DFN1E1 \PLUSETIME180[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[10]_net_1 ));
    DFN1 \CS[16]  (.D(\CS_RNO[16]_net_1 ), .CLK(GLA), .Q(
        \CS[16]_net_1 ));
    XNOR2 fst_lst_pulse_RNO_15 (.A(\necount[3]_net_1 ), .B(
        \NE_NUM[3]_net_1 ), .Y(fst_lst_pulse8_3_i));
    OR2B \timecount_RNO_14[5]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[5]_net_1 ), .Y(\CUTTIME180_TEL_m[5] ));
    OR2B \CS_RNI4H6K[1]  (.A(un1_CS6_39_i_a2_2), .B(N_1343), .Y(
        N_1392_i));
    AOI1B \timecount_RNO_5[9]  (.A(N_1162_i_0), .B(
        \CUTTIME90[9]_net_1 ), .C(\CUTTIME180_m[9] ), .Y(
        timecount_18_iv_9_m1_e_2));
    MX2C \CS_RNO_0[5]  (.A(\CS[5]_net_1 ), .B(\CS[4]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1300));
    DFN1 \CS[14]  (.D(\CS_RNO[14]_net_1 ), .CLK(GLA), .Q(
        \CS[14]_net_1 ));
    MX2 \necount_RNO_0[7]  (.A(\necount1[7] ), .B(\necount[7]_net_1 ), 
        .S(N_1249), .Y(N_518));
    DFN1E0 \CUTTIME180_Tini[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[8]_net_1 ));
    DFN1E0 \OPENTIME[12]  (.D(scaledatain[12]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[12]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E0 \CUTTIME180_TEL[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[6]_net_1 ));
    NOR2B \s_acqnum_1_RNO[0]  (.A(top_code_0_scale_rst), .B(N_348), .Y(
        \s_acqnum_1_RNO[0]_net_1 ));
    DFN1 sw_acq2 (.D(sw_acq2_RNO_3), .CLK(GLA), .Q(
        scalestate_0_sw_acq2));
    DFN1E0 \OPENTIME[2]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[2]_net_1 ));
    DFN1E1 \PLUSETIME90[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[11]_net_1 ));
    OR2B \timecount_RNO_4[5]  (.A(\S_DUMPTIME[5]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[5] ));
    XNOR2 fst_lst_pulse_RNO_8 (.A(\necount[2]_net_1 ), .B(
        \NE_NUM[2]_net_1 ), .Y(fst_lst_pulse8_2_i));
    NOR3C \timecount_RNO_0[5]  (.A(\timecount_18_iv_2[5] ), .B(
        \S_DUMPTIME_m[5] ), .C(\timecount_18_iv_5[5] ), .Y(
        \timecount_18_iv_8[5] ));
    NOR2B \s_acqnum_1_RNO[3]  (.A(top_code_0_scale_rst), .B(N_351), .Y(
        \s_acqnum_1_RNO[3]_net_1 ));
    OR3C \timecount_RNO_3[8]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[8]_net_1 ), .Y(
        \OPENTIME_TEL_m[8] ));
    DFN1E1 \PLUSETIME90[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[5]_net_1 ));
    MX2C \strippluse_RNO_2[9]  (.A(\STRIPNUM90_NUM[9]_net_1 ), .B(
        \STRIPNUM180_NUM[9]_net_1 ), .S(\NS[8] ), .Y(N_245));
    OR2B \timecount_RNO_4[17]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[17]_net_1 ), .Y(\CUTTIME180_m[17] ));
    OR3C \timecount_RNO_6[2]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[2]_net_1 ), .Y(
        \OPENTIME_TEL_m[2] ));
    MX2 \s_acqnum_1_RNO_2[8]  (.A(\ACQ90_NUM[8]_net_1 ), .B(
        \ACQ180_NUM[8]_net_1 ), .S(\NS_0[8] ), .Y(N_272));
    OR2B \timecount_RNO_13[6]  (.A(\S_DUMPTIME[6]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[6] ));
    AOI1B \timecount_RNO_6[10]  (.A(\PLUSETIME180[10]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[10] ), .Y(
        \timecount_18_iv_1[10] ));
    NOR3A DUMPTIME_1_sqmuxa_0_a2 (.A(N_57), .B(N_58), .C(
        scalechoice[0]), .Y(DUMPTIME_1_sqmuxa));
    NOR3C \timecount_RNO_2[8]  (.A(\timecount_18_iv_2[8] ), .B(
        \S_DUMPTIME_m[8] ), .C(\timecount_18_iv_5[8] ), .Y(
        \timecount_18_iv_8[8] ));
    MX2C \CS_RNO_0[19]  (.A(\CS[19]_net_1 ), .B(\CS[3]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1312));
    OR2B \timecount_RNO_8[8]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[8]_net_1 ), .Y(\CUTTIME180_m[8] ));
    AOI1B \timecount_RNO_11[9]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[9]_net_1 ), .C(\CUTTIME180_TEL_m[9] ), .Y(
        timecount_18_iv_9_m1_e_3));
    DFN1E1 \ACQTIME[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[11]_net_1 ));
    XNOR2 M_pulse_RNO_12 (.A(\necount[7]_net_1 ), .B(\M_NUM[7]_net_1 ), 
        .Y(M_pulse8_7_i));
    DFN1 s_acq180 (.D(s_acq180_RNO_net_1), .CLK(GLA), .Q(s_acq180_c));
    DFN1E0 \CUTTIME90[17]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[17]_net_1 ));
    MX2 \s_acqnum_1_RNO_2[3]  (.A(\ACQ90_NUM[3]_net_1 ), .B(
        \ACQ180_NUM[3]_net_1 ), .S(\NS_0[8] ), .Y(N_267));
    DFN1E0 \OPENTIME[7]  (.D(scaledatain[7]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[7]_net_1 ));
    DFN1E1 \ACQECHO_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[6]_net_1 ));
    DFN1E1 \ACQ90_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[9]_net_1 ));
    MX2C \strippluse_RNO_2[5]  (.A(\STRIPNUM90_NUM[5]_net_1 ), .B(
        \STRIPNUM180_NUM[5]_net_1 ), .S(\NS[8] ), .Y(N_241));
    NOR2A \CS_RNO[13]  (.A(top_code_0_scale_rst), .B(N_1307), .Y(
        \CS_RNO[13]_net_1 ));
    OR2B \timecount_RNO_10[7]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[7]_net_1 ), .Y(\CUTTIME180_Tini_m[7] ));
    DFN1E0 \CUTTIME180[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[15]_net_1 ));
    DFN1 \strippluse[7]  (.D(\strippluse_RNO[7]_net_1 ), .CLK(GLA), .Q(
        strippluse[7]));
    OR3C \timecount_RNO[19]  (.A(\timecount_18_0_iv_1[19] ), .B(
        \timecount_18_0_iv_0[19] ), .C(\timecount_18_0_iv_2[19] ), .Y(
        \timecount_18[19] ));
    DFN1E1 \PLUSETIME180[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[7]_net_1 ));
    DFN1E1 \NE_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[2]_net_1 ));
    DFN1E0 \CUTTIME90[8]  (.D(scaledatain[8]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[8]_net_1 ));
    AOI1B \timecount_RNO_5[4]  (.A(N_1162_i_0), .B(
        \CUTTIME90[4]_net_1 ), .C(\CUTTIME180_m[4] ), .Y(
        \timecount_18_iv_2[4] ));
    DFN1E0 \CUTTIME180[4]  (.D(scaledatain[4]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[4]_net_1 ));
    DFN1E1 \ACQ180_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[6]_net_1 ));
    NOR2B long_opentime_RNO (.A(top_code_0_scale_rst), .B(N_525), .Y(
        long_opentime_RNO_net_1));
    AO1C pluse_start_RNO_1 (.A(N_1342), .B(N_1346), .C(N_1278), .Y(
        N_1263));
    DFN1E1 \NE_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[1]_net_1 ));
    DFN1E0 \CUTTIME180[9]  (.D(scaledatain[9]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[9]_net_1 ));
    XA1A fst_lst_pulse_RNO_7 (.A(\NE_NUM[8]_net_1 ), .B(
        \necount[8]_net_1 ), .C(fst_lst_pulse8_4_i), .Y(
        fst_lst_pulse8_NE_3));
    NOR2B \s_acqnum_1_RNO[8]  (.A(top_code_0_scale_rst), .B(N_356), .Y(
        \s_acqnum_1_RNO[8]_net_1 ));
    MX2 reset_out_RNO_0 (.A(N_1323), .B(net_45), .S(N_1245), .Y(N_343));
    NOR3C STRIPNUM90_NUM_1_sqmuxa_0_a2 (.A(N_57), .B(scalechoice[3]), 
        .C(ACQ180_NUM_1_sqmuxa_1), .Y(STRIPNUM90_NUM_1_sqmuxa));
    OR2B \timecount_RNO_13[4]  (.A(\PLUSETIME90[4]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[4] ));
    NOR2B load_out_RNO (.A(top_code_0_scale_rst), .B(N_501), .Y(
        load_out_RNO_net_1));
    DFN1E0 \CUTTIME90[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[14]_net_1 ));
    DFN1E1 \DUMPTIME[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[9]_net_1 ));
    OAI1 \CS_RNO_0[8]  (.A(\CS[8]_net_1 ), .B(
        timer_top_0_clk_en_scale_0), .C(top_code_0_scale_rst), .Y(
        \CS_srsts_i_0[8] ));
    NOR2A \CS_RNO[4]  (.A(top_code_0_scale_rst), .B(N_1299), .Y(
        \CS_RNO_3[4] ));
    DFN1 \CS_i[0]  (.D(\CS_i_RNO_1[0] ), .CLK(GLA), .Q(\CS_i[0]_net_1 )
        );
    MX2 \necount_RNO_0[4]  (.A(\necount1[4] ), .B(\necount[4]_net_1 ), 
        .S(N_1249), .Y(N_515));
    AOI1B \timecount_RNO_5[11]  (.A(\PLUSETIME180[11]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[11] ), .Y(
        \timecount_18_iv_1[11] ));
    NOR2B \CS_RNIUQN4[19]  (.A(top_code_0_scale_rst), .B(
        \CS[19]_net_1 ), .Y(N_1160_i_0));
    DFN1E1 \S_DUMPTIME[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[0]_net_1 ));
    NOR2B \strippluse_RNO[3]  (.A(top_code_0_scale_rst), .B(N_363), .Y(
        \strippluse_RNO[3]_net_1 ));
    NOR2B \necount_RNO[10]  (.A(top_code_0_scale_rst), .B(N_521), .Y(
        \necount_RNO[10]_net_1 ));
    NOR2B \s_acqnum_1_RNO[11]  (.A(top_code_0_scale_rst), .B(N_359), 
        .Y(\s_acqnum_1_RNO[11]_net_1 ));
    DFN1 dds_conf (.D(dds_conf_RNO_1_net_1), .CLK(GLA), .Q(
        scalestate_0_dds_conf));
    DFN1E1 \S_DUMPTIME[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[3]_net_1 ));
    MX2 dump_start_RNO_0 (.A(N_1349), .B(scalestate_0_dump_start), .S(
        N_1251), .Y(N_504));
    MX2C \CS_RNO_0[9]  (.A(\CS[9]_net_1 ), .B(\CS[8]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1303));
    OR2B \timecount_RNO_4[15]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[15]_net_1 ), .Y(\CUTTIME180_TEL_m[15] ));
    MX2 \strippluse_RNO_0[2]  (.A(\strippluse_6[2] ), .B(strippluse[2])
        , .S(un1_CS6_28), .Y(N_362));
    OAI1 \CS_RNITE8C[6]  (.A(\CS[6]_net_1 ), .B(timecount_11_sqmuxa_0), 
        .C(top_code_0_scale_rst), .Y(un1_timecount_5_sqmuxa_3));
    DFN1E0 \CUTTIME180_Tini[20]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[20]_net_1 ));
    AOI1B \timecount_RNO_8[6]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[6]_net_1 ), .C(\OPENTIME_TEL_m[6] ), .Y(
        \timecount_18_iv_4[6] ));
    OR2A \CS_RNII9261[5]  (.A(un1_CS_34_i_a3_0), .B(N_1347), .Y(N_1319)
        );
    MX2C \CS_RNO_0[17]  (.A(\CS[17]_net_1 ), .B(\CS[16]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1311));
    OR3C \timecount_RNO_9[9]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[9]_net_1 ), .Y(
        \OPENTIME_TEL_m[9] ));
    AOI1B \timecount_RNO_13[1]  (.A(N_1162_i_0), .B(
        \CUTTIME90[1]_net_1 ), .C(\CUTTIME180_m[1] ), .Y(
        \timecount_18_iv_10_2[1] ));
    DFN1E1 \PLUSETIME90[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[1]_net_1 ));
    DFN1 \necount[7]  (.D(\necount_RNO[7]_net_1 ), .CLK(GLA), .Q(
        \necount[7]_net_1 ));
    OR2A fst_lst_pulse_RNO (.A(top_code_0_scale_rst), .B(N_523), .Y(
        fst_lst_pulse_RNO_net_1));
    OR3C \timecount_RNO_4[1]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[1]_net_1 ), .Y(
        \OPENTIME_TEL_m[1] ));
    OR2A CS6_0_o2 (.A(top_code_0_scale_rst), .B(
        timer_top_0_clk_en_scale), .Y(N_1278));
    NOR2B off_test_RNO (.A(top_code_0_scale_rst), .B(N_507), .Y(
        off_test_RNO_0_net_1));
    DFN1E1 \timecount[3]  (.D(timecount_18_iv_3_N_2_i_0), .CLK(GLA), 
        .E(un1_CS6_33), .Q(timecount[3]));
    DFN1E0 \OPENTIME_TEL[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[11]_net_1 ));
    DFN1 \strippluse[0]  (.D(\strippluse_RNO[0]_net_1 ), .CLK(GLA), .Q(
        strippluse[0]));
    OR2B \timecount_RNO_4[2]  (.A(\S_DUMPTIME[2]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[2] ));
    NOR2B \strippluse_RNO[0]  (.A(top_code_0_scale_rst), .B(N_360), .Y(
        \strippluse_RNO[0]_net_1 ));
    DFN1E1 \ACQTIME[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[10]_net_1 ));
    AOI1B \timecount_RNO_1[13]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[13]_net_1 ), .C(\CUTTIME180_TEL_m[13] ), .Y(
        \timecount_18_iv_3[13] ));
    OR2B \timecount_RNO_3[17]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[17]_net_1 ), .Y(\CUTTIME180_TEL_m[17] ));
    DFN1E1 \PLUSETIME90[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[3]_net_1 ));
    OR2A intertodsp_RNO_3 (.A(\CS[10]_net_1 ), .B(fst_lst_pulse_net_1), 
        .Y(intertodsp_1_sqmuxa));
    OR2B \timecount_RNO_4[14]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[14]_net_1 ), .Y(\CUTTIME180_TEL_m[14] ));
    MX2 \strippluse_RNO_0[3]  (.A(\strippluse_6[3] ), .B(strippluse[3])
        , .S(un1_CS6_28), .Y(N_363));
    MX2 \s_acqnum_1_RNO_1[3]  (.A(N_267), .B(\ACQECHO_NUM[3]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[3] ));
    MX2 intertodsp_RNO_0 (.A(N_1350), .B(calcuinter_c), .S(un1_CS6_10), 
        .Y(N_508));
    DFN1E0 \CUTTIME180_Tini[19]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[19]_net_1 ));
    NOR2B \CS_RNIOUN4[20]  (.A(top_code_0_scale_rst), .B(
        \CS[20]_net_1 ), .Y(N_1156_i_0));
    DFN1E1 \M_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[0]_net_1 ));
    DFN1E1 \DUMPTIME[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[12]_net_1 ));
    AOI1B \timecount_RNO_0[19]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[19]_net_1 ), .C(\CUTTIME180_TEL_m[19] ), .Y(
        \timecount_18_0_iv_1[19] ));
    NOR2B \CS_RNIQPOA[6]  (.A(top_code_0_scale_rst), .B(\CS[6]_net_1 ), 
        .Y(N_1162_i_0));
    NOR2B M_pulse_RNO (.A(top_code_0_scale_rst), .B(N_527), .Y(
        M_pulse_RNO_net_1));
    DFN1E1 \ACQ90_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[4]_net_1 ));
    AOI1B \timecount_RNO_3[3]  (.A(N_1162_i_0), .B(
        \CUTTIME90[3]_net_1 ), .C(\CUTTIME180_m[3] ), .Y(
        timecount_18_iv_3_m1_e_2));
    OR3C \timecount_RNO_9[4]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[4]_net_1 ), .Y(
        \OPENTIME_TEL_m[4] ));
    AOI1B \timecount_RNO_0[0]  (.A(\S_DUMPTIME[0]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_2[0] ), .Y(
        \timecount_18_iv_6[0] ));
    AND2 \CS_RNI8TMD[18]  (.A(un1_CS6_39_i_a2_1), .B(un1_CS6_39_i_a2_0)
        , .Y(un1_CS6_39_i_a2_2));
    OR3C \timecount_RNO_6[3]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[3]_net_1 ), .Y(
        \OPENTIME_TEL_m[3] ));
    NOR2B \CS_RNIK30D[5]  (.A(N_1346), .B(N_1349), .Y(un1_CS_34_i_a3_0)
        );
    DFN1 \CS[8]  (.D(\CS_RNO_1[8] ), .CLK(GLA), .Q(\CS[8]_net_1 ));
    OR3C \timecount_RNO_5[10]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[10]_net_1 ), .Y(
        \ACQTIME_m[10] ));
    DFN1E0 \CUTTIME180_Tini[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[2]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[0]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[11]_net_1 ));
    DFN1E1 \ACQECHO_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[2]_net_1 ));
    DFN1E1 \timecount[18]  (.D(\timecount_18[18] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[18]));
    MX2 \necount_RNO_0[8]  (.A(\necount1[8] ), .B(\necount[8]_net_1 ), 
        .S(N_1249), .Y(N_519));
    AOI1B \timecount_RNO_1[18]  (.A(N_1162_i_0), .B(
        \CUTTIME90[18]_net_1 ), .C(\CUTTIME180_m[18] ), .Y(
        \timecount_18_0_iv_0[18] ));
    DFN1 \CS[9]  (.D(\CS_RNO_1[9] ), .CLK(GLA), .Q(\CS[9]_net_1 ));
    NOR2B \s_acqnum_1_RNO[2]  (.A(top_code_0_scale_rst), .B(N_350), .Y(
        \s_acqnum_1_RNO[2]_net_1 ));
    NOR2B soft_d_RNO (.A(top_code_0_scale_rst), .B(N_346), .Y(
        soft_d_RNO_2));
    OR3C fst_lst_pulse_RNIJEBD1 (.A(N_1395), .B(sw_acq1_1_sqmuxa), .C(
        N_1278), .Y(un1_CS6_34));
    DFN1E1 \ACQ90_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[6]_net_1 ));
    MX2C \strippluse_RNO_2[1]  (.A(\STRIPNUM90_NUM[1]_net_1 ), .B(
        \STRIPNUM180_NUM[1]_net_1 ), .S(\NS[8] ), .Y(N_237));
    DFN1E1 \PLUSETIME180[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[15]_net_1 ));
    DFN1E1 \timecount[4]  (.D(\timecount_18[4] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[4]));
    DFN1E1 \S_DUMPTIME[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[6]_net_1 ));
    NOR3C \timecount_RNO_1[5]  (.A(\OPENTIME_TEL_m[5] ), .B(
        \CUTTIME180_Tini_m[5] ), .C(\timecount_18_iv_3[5] ), .Y(
        \timecount_18_iv_7[5] ));
    NOR2A ACQ180_NUM_1_sqmuxa_0_a2 (.A(ACQ180_NUM_1_sqmuxa_1), .B(N_63)
        , .Y(ACQ180_NUM_1_sqmuxa));
    DFN1E0 \CUTTIME180[7]  (.D(scaledatain[7]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[7]_net_1 ));
    NOR3C \timecount_RNO_3[9]  (.A(\DUMPTIME_m[9] ), .B(\ACQTIME_m[9] )
        , .C(timecount_18_iv_9_m1_e_1), .Y(timecount_18_iv_9_m1_e_5));
    OR2B \CS_RNI7897[16]  (.A(N_1278), .B(\CS[16]_net_1 ), .Y(N_1255));
    NOR2B pn_out_RNO (.A(top_code_0_scale_rst), .B(N_372), .Y(
        pn_out_RNO_net_1));
    DFN1E1 \PLUSETIME180[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[2]_net_1 ));
    OR3C \timecount_RNO[1]  (.A(\timecount_RNO_0[1]_net_1 ), .B(
        \timecount_18_iv_10_7[1] ), .C(\timecount_18_iv_10_8[1] ), .Y(
        \timecount_18[1] ));
    MX2 \s_acqnum_1_RNO_2[6]  (.A(\ACQ90_NUM[6]_net_1 ), .B(
        \ACQ180_NUM[6]_net_1 ), .S(\NS_0[8] ), .Y(N_270));
    DFN1E1 \STRIPNUM90_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[11]_net_1 ));
    DFN1E1 \DUMPTIME[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[0]_net_1 ));
    MX2 \strippluse_RNO_0[10]  (.A(\strippluse_6[10] ), .B(
        strippluse[10]), .S(un1_CS6_28), .Y(N_370));
    NOR3C \timecount_RNO_5[6]  (.A(\CUTTIME180_m[6] ), .B(
        \CUTTIME90_m[6] ), .C(\S_DUMPTIME_m[6] ), .Y(
        \timecount_18_iv_6[6] ));
    OR3C \timecount_RNO_3[15]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[15]_net_1 ), .Y(
        \OPENTIME_TEL_m[15] ));
    NOR2B \CS_RNI02AS[14]  (.A(timer_top_0_clk_en_scale_0), .B(N_1395), 
        .Y(N_1340));
    OR3C \timecount_RNO_9[11]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[11]_net_1 ), .Y(
        \ACQTIME_m[11] ));
    AOI1B \timecount_RNO_2[9]  (.A(\S_DUMPTIME[9]_net_1 ), .B(
        N_1188_i_0), .C(timecount_18_iv_9_m1_e_2), .Y(
        timecount_18_iv_9_m1_e_6));
    DFN1E1 \S_DUMPTIME[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[11]_net_1 ));
    DFN1E0 \OPENTIME_TEL[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[2]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[14]_net_1 ));
    OR3C \timecount_RNO[5]  (.A(\timecount_18_iv_8[5] ), .B(
        \timecount_18_iv_7[5] ), .C(\timecount_RNO_2[5]_net_1 ), .Y(
        \timecount_18[5] ));
    XNOR2 fst_lst_pulse_RNO_11 (.A(\necount[9]_net_1 ), .B(
        \NE_NUM[9]_net_1 ), .Y(fst_lst_pulse8_9_i));
    AOI1B \timecount_RNO_2[17]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[17]_net_1 ), .C(\OPENTIME_TEL_m[17] ), .Y(
        \timecount_18_0_iv_2[17] ));
    DFN1 necount_LE_NE (.D(necount_LE_NE_RNO_net_1), .CLK(GLA), .Q(
        necount_LE_NE_net_1));
    AO1C pn_out_RNO_2 (.A(\NS[8] ), .B(\CS_i[0]_net_1 ), .C(N_1278), 
        .Y(N_1247));
    NOR2B ACQ180_NUM_1_sqmuxa_0_a2_1 (.A(scalechoice[2]), .B(
        scalechoice[0]), .Y(ACQ180_NUM_1_sqmuxa_1));
    DFN1E0 \CUTTIME180_Tini[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[7]_net_1 ));
    DFN1E1 \ACQTIME[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[7]_net_1 ));
    OA1A dumpoff_ctr_RNO (.A(N_1276), .B(scalestate_0_dumpoff_ctr), .C(
        top_code_0_scale_rst), .Y(dumpoff_ctr_RNO_3));
    MX2 \strippluse_RNO_0[1]  (.A(\strippluse_6[1] ), .B(strippluse[1])
        , .S(un1_CS6_28), .Y(N_361));
    DFN1E1 \S_DUMPTIME[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[7]_net_1 ));
    NOR2B \strippluse_RNO[9]  (.A(top_code_0_scale_rst), .B(N_369), .Y(
        \strippluse_RNO[9]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[15]_net_1 ));
    OR2B \timecount_RNO_14[2]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[2]_net_1 ), .Y(\CUTTIME180_TEL_m[2] ));
    MX2 \strippluse_RNO_0[7]  (.A(\strippluse_6[7] ), .B(strippluse[7])
        , .S(un1_CS6_28), .Y(N_367));
    MX2C \strippluse_RNO_2[2]  (.A(\STRIPNUM90_NUM[2]_net_1 ), .B(
        \STRIPNUM180_NUM[2]_net_1 ), .S(\NS[8] ), .Y(N_238));
    NOR3C ACQTIME_1_sqmuxa_0_a2 (.A(N_57), .B(scalechoice[3]), .C(
        ACQTIME_1_sqmuxa_0_a2_0_net_1), .Y(ACQTIME_1_sqmuxa));
    DFN1E1 \ACQ180_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[9]_net_1 ));
    OR2B \timecount_RNO_12[13]  (.A(\PLUSETIME90[13]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[13] ));
    DFN1E1 \ACQ90_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[0]_net_1 ));
    OR3C \timecount_RNO_3[14]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[14]_net_1 ), .Y(
        \OPENTIME_TEL_m[14] ));
    NOR2A ACQ90_NUM_1_sqmuxa_0_a2_1 (.A(scalechoice[2]), .B(
        scalechoice[0]), .Y(ACQ90_NUM_1_sqmuxa_1));
    NOR3C \timecount_RNO_2[1]  (.A(\timecount_18_iv_10_1[1] ), .B(
        \timecount_18_iv_10_0[1] ), .C(\timecount_18_iv_10_6[1] ), .Y(
        \timecount_18_iv_10_8[1] ));
    DFN1E0 \CUTTIME180_TEL[17]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[17]_net_1 ));
    OR2A rt_sw_RNO_1 (.A(N_1349), .B(N_1348), .Y(N_1318));
    OR2B long_opentime_RNO_1 (.A(timer_top_0_clk_en_scale_0), .B(
        \CS[8]_net_1 ), .Y(N_1267));
    DFN1 \s_acqnum_1[10]  (.D(\s_acqnum_1_RNO[10]_net_1 ), .CLK(GLA), 
        .Q(s_acqnum_1[10]));
    DFN1E1 \NE_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[10]_net_1 ));
    DFN1 reset_out (.D(reset_out_RNO_1_net_1), .CLK(GLA), .Q(net_45));
    DFN1E1 \STRIPNUM180_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[1]_net_1 ));
    NOR3C \timecount_RNO_5[2]  (.A(\DUMPTIME_m[2] ), .B(\ACQTIME_m[2] )
        , .C(\timecount_18_iv_1[2] ), .Y(\timecount_18_iv_5[2] ));
    DFN1E1 \ACQ90_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[5]_net_1 ));
    OR3 OPENTIME_201_e (.A(N_63), .B(scalechoice[2]), .C(
        scalechoice[0]), .Y(N_1436_i));
    OR2B \timecount_RNO_10[15]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[15]_net_1 ), .Y(\CUTTIME180_m[15] ));
    DFN1E1 \PLUSETIME180[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[6]_net_1 ));
    XNOR2 M_pulse_RNO_6 (.A(\necount[5]_net_1 ), .B(\M_NUM[5]_net_1 ), 
        .Y(M_pulse8_5_i));
    DFN1E1 \M_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[6]_net_1 ));
    NOR2B \necount_RNO[4]  (.A(top_code_0_scale_rst), .B(N_515), .Y(
        \necount_RNO[4]_net_1 ));
    AOI1B \timecount_RNO_1[8]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[8]_net_1 ), .C(\CUTTIME180_TEL_m[8] ), .Y(
        \timecount_18_iv_3[8] ));
    DFN1E1 \M_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[7]_net_1 ));
    OR2B \timecount_RNO_11[15]  (.A(N_1162_i_0), .B(
        \CUTTIME90[15]_net_1 ), .Y(\CUTTIME90_m[15] ));
    OR2B \timecount_RNO_8[12]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[12]_net_1 ), .Y(\CUTTIME180_Tini_m[12] ));
    OR3B \timecount_RNO_2[3]  (.A(N_1343), .B(top_code_0_scale_rst), 
        .C(\CS_RNITMND1[6]_net_1 ), .Y(\timecount_RNO_2[3]_net_1 ));
    MX2C \strippluse_RNO_2[10]  (.A(\STRIPNUM90_NUM[10]_net_1 ), .B(
        \STRIPNUM180_NUM[10]_net_1 ), .S(\NS_0[8] ), .Y(N_246));
    NOR2B reset_out_RNO (.A(top_code_0_scale_rst), .B(N_343), .Y(
        reset_out_RNO_1_net_1));
    AOI1B \timecount_RNO_6[0]  (.A(\PLUSETIME180[0]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[0] ), .Y(\timecount_18_iv_1[0] )
        );
    XNOR2 M_pulse_RNO_5 (.A(\necount[6]_net_1 ), .B(\M_NUM[6]_net_1 ), 
        .Y(M_pulse8_6_i));
    DFN1 \strippluse[3]  (.D(\strippluse_RNO[3]_net_1 ), .CLK(GLA), .Q(
        strippluse[3]));
    DFN1E1 \NE_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[9]_net_1 ));
    MX2 \necount_RNO_0[6]  (.A(\necount1[6] ), .B(\necount[6]_net_1 ), 
        .S(N_1249), .Y(N_517));
    MX2C \strippluse_RNO_2[8]  (.A(\STRIPNUM90_NUM[8]_net_1 ), .B(
        \STRIPNUM180_NUM[8]_net_1 ), .S(\NS[8] ), .Y(N_244));
    NOR3C \timecount_RNO_0[3]  (.A(timecount_18_iv_3_m1_e_2), .B(
        \S_DUMPTIME_m[3] ), .C(timecount_18_iv_3_m1_e_5), .Y(
        timecount_18_iv_3_m1_e_8));
    AO1C off_test_RNO_1 (.A(N_1344), .B(N_1346), .C(N_1278), .Y(N_1257)
        );
    DFN1E0 \OPENTIME_TEL[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[14]_net_1 ));
    AOI1B \timecount_RNO_9[10]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[10]_net_1 ), .C(\CUTTIME180_TEL_m[10] ), .Y(
        \timecount_18_iv_3[10] ));
    DFN1 \necount[11]  (.D(\necount_RNO[11]_net_1 ), .CLK(GLA), .Q(
        \necount[11]_net_1 ));
    OR3C \timecount_RNO[3]  (.A(timecount_18_iv_3_m1_e_8), .B(
        timecount_18_iv_3_m1_e_7), .C(\timecount_RNO_2[3]_net_1 ), .Y(
        timecount_18_iv_3_N_2_i_0));
    OR3A \timecount_RNO_2[6]  (.A(top_code_0_scale_rst), .B(N_1347), 
        .C(\CS_RNITMND1[6]_net_1 ), .Y(\timecount_cnst_m[6] ));
    NOR2B M_pulse_RNI9S06 (.A(timecount_16_sqmuxa_1), .B(
        top_code_0_scale_rst), .Y(timecount_16_sqmuxa));
    NOR3C \timecount_RNO_2[15]  (.A(\timecount_18_iv_1[15] ), .B(
        \timecount_18_iv_0[15] ), .C(\timecount_18_iv_6[15] ), .Y(
        \timecount_18_iv_8[15] ));
    DFN1E0 \CUTTIME180[19]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1428), 
        .Q(\CUTTIME180[19]_net_1 ));
    MX2 \s_acqnum_1_RNO_0[5]  (.A(\s_acqnum_7[5] ), .B(s_acqnum_1[5]), 
        .S(un1_CS6_28), .Y(N_353));
    AOI1B \timecount_RNO_0[12]  (.A(\S_DUMPTIME[12]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_2[12] ), .Y(
        \timecount_18_iv_6[12] ));
    DFN1E0 \CUTTIME90[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[13]_net_1 ));
    DFN1E0 \OPENTIME[3]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[3]_net_1 ));
    XNOR2 \necount_RNO_0[0]  (.A(N_1249), .B(\necount[0]_net_1 ), .Y(
        N_511));
    NOR3C M_pulse_RNO_1 (.A(M_pulse8_NE_7), .B(M_pulse8_NE_6), .C(
        M_pulse8_NE_8), .Y(M_pulse8_NE_i_0));
    OR2B \timecount_RNO_4[16]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[16]_net_1 ), .Y(\CUTTIME180_m[16] ));
    NOR3C \timecount_RNO_2[0]  (.A(\OPENTIME_TEL_m[0] ), .B(
        \CUTTIME180_Tini_m[0] ), .C(\timecount_18_iv_3[0] ), .Y(
        \timecount_18_iv_7[0] ));
    DFN1E1 \ACQ90_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[1]_net_1 ));
    MX2 \s_acqnum_1_RNO_1[4]  (.A(N_268), .B(\ACQECHO_NUM[4]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[4] ));
    NOR3C \timecount_RNO_7[15]  (.A(\CUTTIME180_m[15] ), .B(
        \CUTTIME90_m[15] ), .C(\S_DUMPTIME_m[15] ), .Y(
        \timecount_18_iv_6[15] ));
    OR3B CUTTIME90_221_e (.A(N_59), .B(N_62), .C(scalechoice[0]), .Y(
        N_1476_i));
    DFN1E1 \ACQECHO_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[5]_net_1 ));
    DFN1E1 \ACQTIME[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[12]_net_1 ));
    OR2B \timecount_RNO_8[0]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[0]_net_1 ), .Y(\CUTTIME180_Tini_m[0] ));
    DFN1E0 \CUTTIME90[0]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[0]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[4]_net_1 ));
    DFN1E0 \OPENTIME[14]  (.D(scaledatain[14]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[14]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[7]_net_1 ));
    NOR3C \timecount_RNO_5[3]  (.A(\DUMPTIME_m[3] ), .B(\ACQTIME_m[3] )
        , .C(timecount_18_iv_3_m1_e_1), .Y(timecount_18_iv_3_m1_e_5));
    DFN1E1 \timecount[5]  (.D(\timecount_18[5] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[5]));
    OR2B \timecount_RNO_12[14]  (.A(\S_DUMPTIME[14]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[14] ));
    DFN1 \strippluse[5]  (.D(\strippluse_RNO[5]_net_1 ), .CLK(GLA), .Q(
        strippluse[5]));
    MX2C \CS_RNO_0[7]  (.A(\CS[7]_net_1 ), .B(\CS[6]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1302));
    DFN1E1 \S_DUMPTIME[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[1]_net_1 ));
    DFN1E1 \STRIPNUM90_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[1]_net_1 ));
    NOR2 ACQTIME_1_sqmuxa_0_a2_0 (.A(scalechoice[2]), .B(
        scalechoice[0]), .Y(ACQTIME_1_sqmuxa_0_a2_0_net_1));
    DFN1E0 \CUTTIME180_Tini[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[5]_net_1 ));
    NOR2B \s_acqnum_1_RNO[9]  (.A(top_code_0_scale_rst), .B(N_357), .Y(
        \s_acqnum_1_RNO[9]_net_1 ));
    NOR2 \strippluse_RNO_1[4]  (.A(N_240), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[4] ));
    OR3C \timecount_RNO_12[1]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[1]_net_1 ), .Y(
        \ACQTIME_m[1] ));
    MX2C \CS_RNO_0[20]  (.A(\CS[20]_net_1 ), .B(\CS[9]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1313));
    MX2 \necount_RNO_0[10]  (.A(\necount1[10] ), .B(
        \necount[10]_net_1 ), .S(N_1249), .Y(N_521));
    XNOR2 M_pulse_RNO_16 (.A(\necount[10]_net_1 ), .B(
        \M_NUM[10]_net_1 ), .Y(M_pulse8_10_i));
    DFN1E0 \CUTTIME180[17]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1428), 
        .Q(\CUTTIME180[17]_net_1 ));
    DFN1 \CS[7]  (.D(\CS_RNO_3[7] ), .CLK(GLA), .Q(\CS[7]_net_1 ));
    MX2C \CS_RNO_0[10]  (.A(\CS[10]_net_1 ), .B(\CS[20]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1304));
    MX2 dump_sustain_ctrl_RNO_0 (.A(\CS_0[11]_net_1 ), .B(
        scalestate_0_dump_sustain_ctrl), .S(N_1243), .Y(N_526));
    OR3C \timecount_RNO_5[19]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[19]_net_1 ), .Y(
        \OPENTIME_TEL_m[19] ));
    NOR3C \timecount_RNO_2[14]  (.A(\timecount_18_iv_1[14] ), .B(
        \timecount_18_iv_0[14] ), .C(\timecount_18_iv_6[14] ), .Y(
        \timecount_18_iv_8[14] ));
    NOR3C \timecount_RNO_7[14]  (.A(\CUTTIME180_m[14] ), .B(
        \CUTTIME90_m[14] ), .C(\S_DUMPTIME_m[14] ), .Y(
        \timecount_18_iv_6[14] ));
    DFN1 \CS[20]  (.D(\CS_RNO[20]_net_1 ), .CLK(GLA), .Q(
        \CS[20]_net_1 ));
    OR3C OPENTIME_TEL_303_e (.A(N_62), .B(N_64), .C(scalechoice[0]), 
        .Y(N_1640));
    DFN1E1 \ACQTIME[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[0]_net_1 ));
    XNOR2 M_pulse_RNO_9 (.A(\necount[0]_net_1 ), .B(\M_NUM[0]_net_1 ), 
        .Y(M_pulse8_0_i));
    AOI1B \timecount_RNO_6[12]  (.A(\PLUSETIME180[12]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[12] ), .Y(
        \timecount_18_iv_1[12] ));
    DFN1E1 \ACQ90_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[3]_net_1 ));
    OR2B \CS_RNIG7NB[20]  (.A(top_code_0_scale_rst), .B(
        timecount_18_iv_1_m3_e_1), .Y(un1_timecount_5_sqmuxatt_N_6));
    DFN1E0 \CUTTIME180_TEL[19]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[19]_net_1 ));
    DFN1 \CS[6]  (.D(\CS_RNO_3[6] ), .CLK(GLA), .Q(\CS[6]_net_1 ));
    OR2B \timecount_RNO_7[2]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[2]_net_1 ), .Y(\CUTTIME180_Tini_m[2] ));
    DFN1E0 \OPENTIME[15]  (.D(scaledatain[15]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[15]_net_1 ));
    OA1 \CS_i_RNO[0]  (.A(\CS_i[0]_net_1 ), .B(
        timer_top_0_clk_en_scale_0), .C(top_code_0_scale_rst), .Y(
        \CS_i_RNO_1[0] ));
    DFN1E0 \CUTTIME180[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[10]_net_1 ));
    DFN1 \CS[18]  (.D(\CS_RNO[18]_net_1 ), .CLK(GLA), .Q(
        \CS[18]_net_1 ));
    MX2 \strippluse_RNO_0[9]  (.A(\strippluse_6[9] ), .B(strippluse[9])
        , .S(un1_CS6_28), .Y(N_369));
    necount_cmp necount_cmp_0 (.M_NUM({\M_NUM[11]_net_1 , 
        \M_NUM[10]_net_1 , \M_NUM[9]_net_1 , \M_NUM[8]_net_1 , 
        \M_NUM[7]_net_1 , \M_NUM[6]_net_1 , \M_NUM[5]_net_1 , 
        \M_NUM[4]_net_1 , \M_NUM[3]_net_1 , \M_NUM[2]_net_1 , 
        \M_NUM[1]_net_1 , \M_NUM[0]_net_1 }), .necount({
        \necount[11]_net_1 , \necount[10]_net_1 , \necount[9]_net_1 , 
        \necount[8]_net_1 , \necount[7]_net_1 , \necount[6]_net_1 , 
        \necount[5]_net_1 , \necount[4]_net_1 , \necount[3]_net_1 , 
        \necount[2]_net_1 , \necount[1]_net_1 , \necount[0]_net_1 }), 
        .necount_LE_M_1(necount_LE_M_1));
    MX2 \s_acqnum_1_RNO_1[2]  (.A(N_266), .B(\ACQECHO_NUM[2]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[2] ));
    DFN1E1 \timecount[9]  (.D(timecount_18_iv_9_N_2_i_0), .CLK(GLA), 
        .E(un1_CS6_33), .Q(timecount[9]));
    DFN1E0 \CUTTIME180[18]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1428), 
        .Q(\CUTTIME180[18]_net_1 ));
    DFN1E1 \ACQTIME[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[2]_net_1 ));
    NOR3C \timecount_RNO_1[1]  (.A(\OPENTIME_TEL_m[1] ), .B(
        \CUTTIME180_Tini_m[1] ), .C(\timecount_18_iv_10_3[1] ), .Y(
        \timecount_18_iv_10_7[1] ));
    MX2 \s_acqnum_1_RNO_2[7]  (.A(\ACQ90_NUM[7]_net_1 ), .B(
        \ACQ180_NUM[7]_net_1 ), .S(\NS_0[8] ), .Y(N_271));
    DFN1E1 \DUMPTIME[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[15]_net_1 ));
    DFN1 \necount[4]  (.D(\necount_RNO[4]_net_1 ), .CLK(GLA), .Q(
        \necount[4]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[10]_net_1 ));
    DFN1E1 \STRIPNUM90_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[9]_net_1 ));
    DFN1E1 \ACQ90_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[11]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[3]_net_1 ));
    NOR3C ACQECHO_NUM_1_sqmuxa_0_a2 (.A(N_57), .B(scalechoice[3]), .C(
        ACQ90_NUM_1_sqmuxa_1), .Y(ACQECHO_NUM_1_sqmuxa));
    AO1B tetw_pluse_RNO (.A(scalestate_0_tetw_pluse), .B(N_1276), .C(
        top_code_0_scale_rst), .Y(tetw_pluse_RNO_0));
    MX2 \necount_RNO_0[5]  (.A(\necount1[5] ), .B(\necount[5]_net_1 ), 
        .S(N_1249), .Y(N_516));
    MX2 \s_acqnum_1_RNO_1[6]  (.A(N_270), .B(\ACQECHO_NUM[6]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[6] ));
    DFN1E0 \OPENTIME_TEL[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[7]_net_1 ));
    OR3C intertodsp_RNO_1 (.A(N_1322), .B(intertodsp_1_sqmuxa), .C(
        N_1278), .Y(un1_CS6_10));
    XNOR2 fst_lst_pulse_RNO_9 (.A(\necount[0]_net_1 ), .B(
        \NE_NUM[0]_net_1 ), .Y(fst_lst_pulse8_0_i));
    NOR2A un1_PLUSETIME9030_1_i_a2_0 (.A(scalechoice[2]), .B(
        scalechoice[3]), .Y(N_62));
    DFN1E1 \STRIPNUM90_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[10]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[14]_net_1 ));
    NOR2B \necount_RNO[7]  (.A(top_code_0_scale_rst), .B(N_518), .Y(
        \necount_RNO[7]_net_1 ));
    OR3C CUTTIME90_237_e (.A(N_59), .B(N_62), .C(scalechoice[0]), .Y(
        N_1508));
    DFN1E1 \PLUSETIME180[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[12]_net_1 ));
    MX2A sw_acq1_RNO_0 (.A(N_1347), .B(scalestate_0_sw_acq1), .S(
        un1_CS6_34), .Y(N_345));
    NOR2B M_pulse_RNI9S06_0 (.A(timecount_15_sqmuxa_1), .B(
        top_code_0_scale_rst), .Y(timecount_15_sqmuxa));
    DFN1E0 \CUTTIME90[3]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[3]_net_1 ));
    OR2B \timecount_RNO_3[16]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[16]_net_1 ), .Y(\CUTTIME180_TEL_m[16] ));
    DFN1E0 \CUTTIME180_TEL[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[0]_net_1 ));
    DFN1E1 \S_DUMPTIME[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[4]_net_1 ));
    DFN1E1 \timecount[1]  (.D(\timecount_18[1] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[1]));
    DFN1E0 \OPENTIME[0]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[0]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[11]_net_1 ));
    NOR3B M_pulse_RNIVLG1 (.A(M_pulse_net_1), .B(\CS[15]_net_1 ), .C(
        necount_LE_M_net_1), .Y(timecount_15_sqmuxa_1));
    OR2B \timecount_RNO_4[8]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[8]_net_1 ), .Y(\CUTTIME180_TEL_m[8] ));
    MX2 \s_acqnum_1_RNO_2[10]  (.A(\ACQ90_NUM[10]_net_1 ), .B(
        \ACQ180_NUM[10]_net_1 ), .S(\NS[8] ), .Y(N_274));
    DFN1E1 \S_DUMPTIME[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[5]_net_1 ));
    NOR3B \CS_RNO_0[18]  (.A(\CS[17]_net_1 ), .B(
        timer_top_0_clk_en_scale), .C(necount_LE_NE_net_1), .Y(N_1289));
    NOR2B \necount_RNO[5]  (.A(top_code_0_scale_rst), .B(N_516), .Y(
        \necount_RNO[5]_net_1 ));
    DFN1E1 \ACQ180_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[3]_net_1 ));
    NOR3C \timecount_RNO_1[3]  (.A(\OPENTIME_TEL_m[3] ), .B(
        \CUTTIME180_Tini_m[3] ), .C(timecount_18_iv_3_m1_e_3), .Y(
        timecount_18_iv_3_m1_e_7));
    DFN1E1 \ACQECHO_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[4]_net_1 ));
    NOR2B \s_acqnum_1_RNO[4]  (.A(top_code_0_scale_rst), .B(N_352), .Y(
        \s_acqnum_1_RNO[4]_net_1 ));
    DFN1 \CS[15]  (.D(\CS_RNO[15]_net_1 ), .CLK(GLA), .Q(
        \CS[15]_net_1 ));
    OR3C \timecount_RNO_7[9]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[9]_net_1 ), .Y(
        \ACQTIME_m[9] ));
    OR3C \timecount_RNO_7[7]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[7]_net_1 ), .Y(
        \ACQTIME_m[7] ));
    AO1 \CS_RNIVM7D_0[7]  (.A(necount_LE_NE_net_1), .B(\CS[17]_net_1 ), 
        .C(\CS[7]_net_1 ), .Y(\NS_0[8] ));
    AOI1B \timecount_RNO_8[9]  (.A(\PLUSETIME180[9]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[9] ), .Y(
        timecount_18_iv_9_m1_e_1));
    OR2B \timecount_RNO_4[11]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[11]_net_1 ), .Y(\CUTTIME180_TEL_m[11] ));
    DFN1E0 \CUTTIME90[18]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[18]_net_1 ));
    DFN1E1 \S_DUMPTIME[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[13]_net_1 ));
    DFN1 necount_LE_M (.D(necount_LE_M_RNO_net_1), .CLK(GLA), .Q(
        necount_LE_M_net_1));
    MX2 \s_acqnum_1_RNO_0[10]  (.A(\s_acqnum_7[10] ), .B(
        s_acqnum_1[10]), .S(un1_CS6_28), .Y(N_358));
    MX2 pluse_start_RNO_0 (.A(N_1342), .B(scalestate_0_pluse_start), 
        .S(N_1263), .Y(N_506));
    MX2 \s_acqnum_1_RNO_1[7]  (.A(N_271), .B(\ACQECHO_NUM[7]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[7] ));
    NOR2B rt_sw_RNO (.A(top_code_0_scale_rst), .B(N_347), .Y(
        rt_sw_RNO_4));
    DFN1E1 \S_DUMPTIME[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[15]_net_1 ));
    AOI1B \timecount_RNO_4[6]  (.A(N_1185_i_0), .B(\DUMPTIME[6]_net_1 )
        , .C(\ACQTIME_m[6] ), .Y(\timecount_18_iv_0[6] ));
    MX2 \s_acqnum_1_RNO_0[6]  (.A(\s_acqnum_7[6] ), .B(s_acqnum_1[6]), 
        .S(un1_CS6_28), .Y(N_354));
    DFN1E0 \CUTTIME90[1]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[1]_net_1 ));
    OR3C \timecount_RNO_11[3]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[3]_net_1 ), .Y(
        \ACQTIME_m[3] ));
    DFN1E1 \NE_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[5]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[11]_net_1 ));
    OR2 \CS_RNI5RHC[8]  (.A(\CS[9]_net_1 ), .B(\CS[8]_net_1 ), .Y(
        N_1320));
    NOR2B \necount_RNO[9]  (.A(top_code_0_scale_rst), .B(N_520), .Y(
        \necount_RNO[9]_net_1 ));
    OR2B \timecount_RNO_8[13]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[13]_net_1 ), .Y(\CUTTIME180_m[13] ));
    AOI1B \timecount_RNO_6[1]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[1]_net_1 ), .C(\CUTTIME180_TEL_m[1] ), .Y(
        \timecount_18_iv_10_3[1] ));
    OR2B \timecount_RNO_10[10]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[10]_net_1 ), .Y(\CUTTIME180_m[10] ));
    DFN1E1 \ACQECHO_NUM[3]  (.D(scaledatain[3]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[3]_net_1 ));
    DFN1E1 \ACQECHO_NUM[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[1]_net_1 ));
    MX2C \CS_RNO_0[14]  (.A(\CS[14]_net_1 ), .B(\CS[13]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1308));
    DFN1E0 \OPENTIME[18]  (.D(scaledatain[2]), .CLK(GLA), .E(N_1468), 
        .Q(\OPENTIME[18]_net_1 ));
    OR2B \timecount_RNO_11[10]  (.A(\PLUSETIME90[10]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[10] ));
    OR3C \timecount_RNO_5[12]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[12]_net_1 ), .Y(
        \ACQTIME_m[12] ));
    DFN1E0 \OPENTIME_TEL[20]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[20]_net_1 ));
    DFN1 \s_acqnum_1[0]  (.D(\s_acqnum_1_RNO[0]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[0]));
    DFN1 \necount[1]  (.D(\necount_RNO[1]_net_1 ), .CLK(GLA), .Q(
        \necount[1]_net_1 ));
    OR3B CUTTIME180_TEL_259_e (.A(un1_PLUSETIME9030_3_i_a2_0_net_1), 
        .B(scalechoice[0]), .C(N_58), .Y(N_1552));
    AOI1B \timecount_RNO_0[13]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[13]_net_1 ), .C(\OPENTIME_TEL_m[13] ), .Y(
        \timecount_18_iv_4[13] ));
    NOR2B \strippluse_RNO[4]  (.A(top_code_0_scale_rst), .B(N_364), .Y(
        \strippluse_RNO[4]_net_1 ));
    NOR3B \timecount_RNO_9[5]  (.A(N_1343), .B(top_code_0_scale_rst), 
        .C(N_1342), .Y(N_1337));
    AOI1B \timecount_RNO_2[16]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[16]_net_1 ), .C(\OPENTIME_TEL_m[16] ), .Y(
        \timecount_18_0_iv_2[16] ));
    DFN1E1 \ACQECHO_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[9]_net_1 ));
    NOR2B \strippluse_RNO[8]  (.A(top_code_0_scale_rst), .B(N_368), .Y(
        \strippluse_RNO[8]_net_1 ));
    DFN1E1 \timecount[17]  (.D(\timecount_18[17] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[17]));
    DFN1 \s_acqnum_1[1]  (.D(\s_acqnum_1_RNO[1]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[1]));
    DFN1E1 \PLUSETIME180[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[1]_net_1 ));
    DFN1E1 \timecount[7]  (.D(\timecount_18[7] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[7]));
    DFN1 \CS[13]  (.D(\CS_RNO[13]_net_1 ), .CLK(GLA), .Q(
        \CS[13]_net_1 ));
    DFN1E0 \CUTTIME90[9]  (.D(scaledatain[9]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[9]_net_1 ));
    DFN1 \necount[6]  (.D(\necount_RNO[6]_net_1 ), .CLK(GLA), .Q(
        \necount[6]_net_1 ));
    NOR2 \strippluse_RNO_1[3]  (.A(N_239), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[3] ));
    DFN1E1 \ACQTIME[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[4]_net_1 ));
    DFN1 \CS[3]  (.D(\CS_RNO_3[3] ), .CLK(GLA), .Q(\CS[3]_net_1 ));
    AOI1B \timecount_RNO_8[4]  (.A(\PLUSETIME180[4]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[4] ), .Y(\timecount_18_iv_1[4] )
        );
    OR2B \timecount_RNO_10[0]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[0]_net_1 ), .Y(\CUTTIME180_m[0] ));
    DFN1E1 \PLUSETIME90[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[2]_net_1 ));
    NOR2 \strippluse_RNO_1[11]  (.A(N_247), .B(\CS_0[11]_net_1 ), .Y(
        \strippluse_6[11] ));
    DFN1 soft_d (.D(soft_d_RNO_2), .CLK(GLA), .Q(scalestate_0_soft_d));
    DFN1E0 \CUTTIME180_TEL[21]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[21]_net_1 ));
    OR2B \timecount_RNO_11[2]  (.A(N_1185_i_0), .B(\DUMPTIME[2]_net_1 )
        , .Y(\DUMPTIME_m[2] ));
    OR3 \CS_RNIF0HN[1]  (.A(\CS_0[11]_net_1 ), .B(\CS[1]_net_1 ), .C(
        \NS_0[8] ), .Y(N_1179));
    DFN1E1 \ACQ180_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[5]_net_1 ));
    OR2B \timecount_RNO_4[10]  (.A(N_1185_i_0), .B(
        \DUMPTIME[10]_net_1 ), .Y(\DUMPTIME_m[10] ));
    MX2 \strippluse_RNO_0[5]  (.A(\strippluse_6[5] ), .B(strippluse[5])
        , .S(un1_CS6_28), .Y(N_365));
    OR3B OPENTIME_TEL_287_e (.A(N_62), .B(N_64), .C(scalechoice[0]), 
        .Y(N_1608_i));
    MX2C \strippluse_RNO_2[4]  (.A(\STRIPNUM90_NUM[4]_net_1 ), .B(
        \STRIPNUM180_NUM[4]_net_1 ), .S(\NS[8] ), .Y(N_240));
    OR2A \CS_RNIU52P[2]  (.A(N_1345), .B(N_1342), .Y(N_1347));
    DFN1E1 \DUMPTIME[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[11]_net_1 ));
    AOI1B \timecount_RNO_0[18]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[18]_net_1 ), .C(\CUTTIME180_TEL_m[18] ), .Y(
        \timecount_18_0_iv_1[18] ));
    OR3B CUTTIME180_181_e (.A(N_57), .B(N_62), .C(scalechoice[0]), .Y(
        N_1396_i));
    OR2B \timecount_RNO_6[4]  (.A(N_1185_i_0), .B(\DUMPTIME[4]_net_1 ), 
        .Y(\DUMPTIME_m[4] ));
    NOR3C M_pulse_RNO_2 (.A(M_pulse8_6_i), .B(M_pulse8_5_i), .C(
        M_pulse8_NE_3), .Y(M_pulse8_NE_7));
    DFN1 \strippluse[6]  (.D(\strippluse_RNO[6]_net_1 ), .CLK(GLA), .Q(
        strippluse[6]));
    AOI1B \timecount_RNO_3[6]  (.A(\PLUSETIME180[6]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[6] ), .Y(\timecount_18_iv_1[6] )
        );
    MX2 \s_acqnum_1_RNO_1[1]  (.A(N_265), .B(\ACQECHO_NUM[1]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[1] ));
    DFN1E1 \ACQ90_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[8]_net_1 ));
    MX2C \CS_RNO_0[3]  (.A(\CS[3]_net_1 ), .B(\CS[2]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1298));
    OR2B \timecount_RNO_10[5]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[5]_net_1 ), .Y(\CUTTIME180_m[5] ));
    DFN1 off_test (.D(off_test_RNO_0_net_1), .CLK(GLA), .Q(
        scalestate_0_off_test));
    OR3C \timecount_RNO_10[8]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[8]_net_1 ), .Y(
        \ACQTIME_m[8] ));
    DFN1E0 \CUTTIME180_TEL[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[5]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[10]_net_1 ));
    OR2B \timecount_RNO_6[13]  (.A(\S_DUMPTIME[13]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[13] ));
    AOI1B \timecount_RNO_3[0]  (.A(N_1162_i_0), .B(
        \CUTTIME90[0]_net_1 ), .C(\CUTTIME180_m[0] ), .Y(
        \timecount_18_iv_2[0] ));
    OR3C \timecount_RNO[16]  (.A(\timecount_18_0_iv_1[16] ), .B(
        \timecount_18_0_iv_0[16] ), .C(\timecount_18_0_iv_2[16] ), .Y(
        \timecount_18[16] ));
    OR3C \timecount_RNO[15]  (.A(\timecount_18_iv_4[15] ), .B(
        \timecount_18_iv_3[15] ), .C(\timecount_18_iv_8[15] ), .Y(
        \timecount_18[15] ));
    DFN1E1 \STRIPNUM180_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[7]_net_1 ));
    DFN1E0 \CUTTIME180[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[13]_net_1 ));
    NOR2A \CS_RNO[3]  (.A(top_code_0_scale_rst), .B(N_1298), .Y(
        \CS_RNO_3[3] ));
    AOI1B \timecount_RNO_1[17]  (.A(N_1162_i_0), .B(
        \CUTTIME90[17]_net_1 ), .C(\CUTTIME180_m[17] ), .Y(
        \timecount_18_0_iv_0[17] ));
    DFN1 \necount[3]  (.D(\necount_RNO[3]_net_1 ), .CLK(GLA), .Q(
        \necount[3]_net_1 ));
    OR3C \timecount_RNO_3[11]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[11]_net_1 ), .Y(
        \OPENTIME_TEL_m[11] ));
    DFN1E1 \STRIPNUM90_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[4]_net_1 ));
    NOR3C fst_lst_pulse_RNO_3 (.A(fst_lst_pulse8_2_i), .B(
        fst_lst_pulse8_0_i), .C(fst_lst_pulse8_NE_1), .Y(
        fst_lst_pulse8_NE_6));
    OR3C \timecount_RNO_0[1]  (.A(\timecount_RNO_3[1]_net_1 ), .B(
        un1_timecount_5_sqmuxa_3), .C(un1_timecount_5_sqmuxa_5), .Y(
        \timecount_RNO_0[1]_net_1 ));
    DFN1 \necount[10]  (.D(\necount_RNO[10]_net_1 ), .CLK(GLA), .Q(
        \necount[10]_net_1 ));
    DFN1E1 \S_DUMPTIME[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[9]_net_1 ));
    DFN1E0 \OPENTIME[1]  (.D(scaledatain[1]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[1]_net_1 ));
    DFN1 \CS[10]  (.D(\CS_RNO[10]_net_1 ), .CLK(GLA), .Q(
        \CS[10]_net_1 ));
    DFN1 intertodsp (.D(intertodsp_RNO_0_net_1), .CLK(GLA), .Q(
        calcuinter_c));
    OR2B \timecount_RNO_12[6]  (.A(N_1162_i_0), .B(
        \CUTTIME90[6]_net_1 ), .Y(\CUTTIME90_m[6] ));
    DFN1E1 \timecount[8]  (.D(\timecount_18[8] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[8]));
    OR2 s_acq_RNO_2 (.A(\CS[4]_net_1 ), .B(\CS[15]_net_1 ), .Y(
        un1_CS6_17_i_a3_0));
    DFN1E1 \NE_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[8]_net_1 ));
    NOR3A M_pulse_RNIVLG1_0 (.A(\CS[15]_net_1 ), .B(necount_LE_M_net_1)
        , .C(M_pulse_net_1), .Y(timecount_16_sqmuxa_1));
    DFN1E0 \CUTTIME180_TEL[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[12]_net_1 ));
    DFN1E0 \OPENTIME[6]  (.D(scaledatain[6]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[6]_net_1 ));
    DFN1E1 \ACQ90_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[10]_net_1 ));
    NOR2B dds_conf_RNO (.A(top_code_0_scale_rst), .B(N_509), .Y(
        dds_conf_RNO_1_net_1));
    DFN1E1 \NE_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[11]_net_1 ));
    MX2 dds_conf_RNO_0 (.A(N_1347), .B(scalestate_0_dds_conf), .S(
        N_1265), .Y(N_509));
    OR2B \timecount_RNO_12[11]  (.A(\S_DUMPTIME[11]_net_1 ), .B(
        N_1188_i_0), .Y(\S_DUMPTIME_m[11] ));
    MX2 \s_acqnum_1_RNO_0[4]  (.A(\s_acqnum_7[4] ), .B(s_acqnum_1[4]), 
        .S(un1_CS6_28), .Y(N_352));
    OR2B \timecount_RNO_11[0]  (.A(\PLUSETIME90[0]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[0] ));
    NOR2 \CS_RNI59F[18]  (.A(\CS[18]_net_1 ), .B(\CS[17]_net_1 ), .Y(
        un1_CS6_39_i_a2_1));
    DFN1E1 \STRIPNUM180_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[2]_net_1 ));
    DFN1 dump_start (.D(dump_start_RNO_2), .CLK(GLA), .Q(
        scalestate_0_dump_start));
    DFN1E0 \OPENTIME[16]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1468), 
        .Q(\OPENTIME[16]_net_1 ));
    XNOR2 fst_lst_pulse_RNO_12 (.A(\necount[7]_net_1 ), .B(
        \NE_NUM[7]_net_1 ), .Y(fst_lst_pulse8_7_i));
    DFN1 \strippluse[4]  (.D(\strippluse_RNO[4]_net_1 ), .CLK(GLA), .Q(
        strippluse[4]));
    DFN1E0 \CUTTIME180_Tini[17]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[17]_net_1 ));
    DFN1E1 \STRIPNUM90_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[8]_net_1 ));
    DFN1 \necount[5]  (.D(\necount_RNO[5]_net_1 ), .CLK(GLA), .Q(
        \necount[5]_net_1 ));
    AOI1B \timecount_RNO_9[12]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[12]_net_1 ), .C(\CUTTIME180_TEL_m[12] ), .Y(
        \timecount_18_iv_3[12] ));
    DFN1E0 \OPENTIME_TEL[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[8]_net_1 ));
    DFN1E1 \ACQECHO_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[7]_net_1 ));
    AOI1B \timecount_RNO_12[3]  (.A(\PLUSETIME180[3]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[3] ), .Y(
        timecount_18_iv_3_m1_e_1));
    OA1 \CS_RNI5A0B[5]  (.A(\CS[5]_net_1 ), .B(\CS[11]_net_1 ), .C(
        top_code_0_scale_rst), .Y(N_1188_i_0));
    OR3C \timecount_RNO[21]  (.A(\OPENTIME_TEL_m[21] ), .B(
        \CUTTIME180_Tini_m[21] ), .C(\timecount_18_0_iv_0[21] ), .Y(
        \timecount_18[21] ));
    MX2 soft_d_RNO_0 (.A(scalestate_0_soft_d), .B(N_1319), .S(N_1340), 
        .Y(N_346));
    DFN1E0 \CUTTIME90[5]  (.D(scaledatain[5]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[5]_net_1 ));
    DFN1 long_opentime (.D(long_opentime_RNO_net_1), .CLK(GLA), .Q(
        scalestate_0_long_opentime));
    NOR3B PLUSETIME180_1_sqmuxa_0_a2 (.A(scalechoice[0]), .B(N_59), .C(
        N_58), .Y(PLUSETIME180_1_sqmuxa));
    XNOR2 M_pulse_RNO_11 (.A(\necount[9]_net_1 ), .B(\M_NUM[9]_net_1 ), 
        .Y(M_pulse8_9_i));
    AOI1B \timecount_RNO_1[15]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[15]_net_1 ), .C(\CUTTIME180_TEL_m[15] ), .Y(
        \timecount_18_iv_3[15] ));
    DFN1E1 \PLUSETIME90[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[9]_net_1 ));
    MX2 rt_sw_RNO_0 (.A(scalestate_0_rt_sw), .B(N_1318), .S(N_1340), 
        .Y(N_347));
    DFN1E0 \OPENTIME[8]  (.D(scaledatain[8]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[8]_net_1 ));
    AOI1B \timecount_RNO_3[10]  (.A(N_1162_i_0), .B(
        \CUTTIME90[10]_net_1 ), .C(\CUTTIME180_m[10] ), .Y(
        \timecount_18_iv_2[10] ));
    AOI1B \timecount_RNO_2[4]  (.A(\S_DUMPTIME[4]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_2[4] ), .Y(
        \timecount_18_iv_6[4] ));
    MX2 \s_acqnum_1_RNO_2[5]  (.A(\ACQ90_NUM[5]_net_1 ), .B(
        \ACQ180_NUM[5]_net_1 ), .S(\NS_0[8] ), .Y(N_269));
    MX2 long_opentime_RNO_0 (.A(necount_LE_M_net_1), .B(
        scalestate_0_long_opentime), .S(N_1267), .Y(N_525));
    NOR2B \s_acqnum_1_RNO[1]  (.A(top_code_0_scale_rst), .B(N_349), .Y(
        \s_acqnum_1_RNO[1]_net_1 ));
    NOR2 \CS_RNIR3G6[5]  (.A(\CS[11]_net_1 ), .B(\CS[5]_net_1 ), .Y(
        N_1349));
    OR2B \timecount_RNO_12[12]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[12]_net_1 ), .Y(\CUTTIME180_TEL_m[12] ));
    OR3C \timecount_RNO[17]  (.A(\timecount_18_0_iv_1[17] ), .B(
        \timecount_18_0_iv_0[17] ), .C(\timecount_18_0_iv_2[17] ), .Y(
        \timecount_18[17] ));
    NOR3C \timecount_RNO_2[11]  (.A(\timecount_18_iv_1[11] ), .B(
        \timecount_18_iv_0[11] ), .C(\timecount_18_iv_6[11] ), .Y(
        \timecount_18_iv_8[11] ));
    DFN1E0 \OPENTIME[5]  (.D(scaledatain[5]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[5]_net_1 ));
    OR3C \timecount_RNO_9[7]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[7]_net_1 ), .Y(
        \OPENTIME_TEL_m[7] ));
    OR3C \timecount_RNO[11]  (.A(\timecount_18_iv_4[11] ), .B(
        \timecount_18_iv_3[11] ), .C(\timecount_18_iv_8[11] ), .Y(
        \timecount_18[11] ));
    NOR3C \timecount_RNO_7[11]  (.A(\CUTTIME180_m[11] ), .B(
        \CUTTIME90_m[11] ), .C(\S_DUMPTIME_m[11] ), .Y(
        \timecount_18_iv_6[11] ));
    DFN1 \necount[0]  (.D(\necount_RNO[0]_net_1 ), .CLK(GLA), .Q(
        \necount[0]_net_1 ));
    DFN1 \necount[2]  (.D(\necount_RNO[2]_net_1 ), .CLK(GLA), .Q(
        \necount[2]_net_1 ));
    DFN1E0 \CUTTIME180[8]  (.D(scaledatain[8]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[8]_net_1 ));
    NOR2B \s_acqnum_1_RNO[6]  (.A(top_code_0_scale_rst), .B(N_354), .Y(
        \s_acqnum_1_RNO[6]_net_1 ));
    NOR3C NE_NUM_1_sqmuxa_0_a2 (.A(N_57), .B(scalechoice[3]), .C(
        NE_NUM_1_sqmuxa_0_a2_0_net_1), .Y(NE_NUM_1_sqmuxa));
    DFN1 \s_acqnum_1[9]  (.D(\s_acqnum_1_RNO[9]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[9]));
    MX2 \s_acqnum_1_RNO_2[11]  (.A(\ACQ90_NUM[11]_net_1 ), .B(
        \ACQ180_NUM[11]_net_1 ), .S(\NS[8] ), .Y(N_275));
    OR3C \CS_RNITMND1[6]  (.A(un1_timecount_5_sqmuxatt_N_6), .B(
        un1_timecount_5_sqmuxa_3), .C(un1_timecount_5_sqmuxa_5), .Y(
        \CS_RNITMND1[6]_net_1 ));
    OR2B \timecount_RNO_11[6]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[6]_net_1 ), .Y(\CUTTIME180_m[6] ));
    MX2 \necount_RNO_0[3]  (.A(\necount1[3] ), .B(\necount[3]_net_1 ), 
        .S(N_1249), .Y(N_514));
    DFN1E1 \ACQ90_NUM[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[7]_net_1 ));
    necount_inc necount_inc_0 (.necount({\necount[11]_net_1 , 
        \necount[10]_net_1 , \necount[9]_net_1 , \necount[8]_net_1 , 
        \necount[7]_net_1 , \necount[6]_net_1 , \necount[5]_net_1 , 
        \necount[4]_net_1 , \necount[3]_net_1 , \necount[2]_net_1 , 
        \necount[1]_net_1 , \necount[0]_net_1 }), .necount1({
        \necount1[11] , \necount1[10] , \necount1[9] , \necount1[8] , 
        \necount1[7] , \necount1[6] , \necount1[5] , \necount1[4] , 
        \necount1[3] , \necount1[2] , \necount1[1] }));
    AOI1B \timecount_RNO_1[14]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[14]_net_1 ), .C(\CUTTIME180_TEL_m[14] ), .Y(
        \timecount_18_iv_3[14] ));
    DFN1E1 \PLUSETIME90[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[0]_net_1 ));
    OR2B \timecount_RNO_13[9]  (.A(\PLUSETIME90[9]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[9] ));
    NOR2A \CS_RNO[19]  (.A(top_code_0_scale_rst), .B(N_1312), .Y(
        \CS_RNO[19]_net_1 ));
    OR3C \timecount_RNO_12[2]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[2]_net_1 ), .Y(
        \ACQTIME_m[2] ));
    AOI1B \timecount_RNO_5[13]  (.A(N_1162_i_0), .B(
        \CUTTIME90[13]_net_1 ), .C(\CUTTIME180_m[13] ), .Y(
        \timecount_18_iv_2[13] ));
    MX2 \strippluse_RNO_0[8]  (.A(\strippluse_6[8] ), .B(strippluse[8])
        , .S(un1_CS6_28), .Y(N_368));
    DFN1 \necount[8]  (.D(\necount_RNO[8]_net_1 ), .CLK(GLA), .Q(
        \necount[8]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[6]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[13]_net_1 ));
    DFN1 \CS[19]  (.D(\CS_RNO[19]_net_1 ), .CLK(GLA), .Q(
        \CS[19]_net_1 ));
    MX2 \s_acqnum_1_RNO_0[11]  (.A(\s_acqnum_7[11] ), .B(
        s_acqnum_1[11]), .S(un1_CS6_28), .Y(N_359));
    OR2B \timecount_RNO_7[5]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[5]_net_1 ), .Y(\CUTTIME180_Tini_m[5] ));
    DFN1 pn_out (.D(pn_out_RNO_net_1), .CLK(GLA), .Q(
        scalestate_0_pn_out));
    MX2 off_test_RNO_0 (.A(N_1344), .B(scalestate_0_off_test), .S(
        N_1257), .Y(N_507));
    OR2B \timecount_RNO_4[19]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[19]_net_1 ), .Y(\CUTTIME180_m[19] ));
    DFN1 \s_acqnum_1[5]  (.D(\s_acqnum_1_RNO[5]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[5]));
    DFN1E1 \M_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[8]_net_1 ));
    DFN1E1 \PLUSETIME90[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[13]_net_1 ));
    MX2 \necount_RNO_0[1]  (.A(\necount1[1] ), .B(\necount[1]_net_1 ), 
        .S(N_1249), .Y(N_512));
    DFN1 M_pulse (.D(M_pulse_RNO_net_1), .CLK(GLA), .Q(M_pulse_net_1));
    DFN1 \CS[2]  (.D(\CS_RNO_3[2] ), .CLK(GLA), .Q(\CS[2]_net_1 ));
    NOR2B \timecount_RNO_0[9]  (.A(N_1342), .B(top_code_0_scale_rst), 
        .Y(timecount_18_ivtt_9_m1_e_0));
    DFN1E1 \ACQECHO_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[8]_net_1 ));
    AOI1B \timecount_RNO_3[5]  (.A(N_1162_i_0), .B(
        \CUTTIME90[5]_net_1 ), .C(\CUTTIME180_m[5] ), .Y(
        \timecount_18_iv_2[5] ));
    DFN1E0 \OPENTIME_TEL[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[9]_net_1 ));
    AOI1B \timecount_RNO_11[7]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[7]_net_1 ), .C(\CUTTIME180_TEL_m[7] ), .Y(
        \timecount_18_iv_3[7] ));
    DFN1 \s_acqnum_1[3]  (.D(\s_acqnum_1_RNO[3]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[3]));
    DFN1E1 \timecount[11]  (.D(\timecount_18[11] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[11]));
    NOR2B \necount_RNO[1]  (.A(top_code_0_scale_rst), .B(N_512), .Y(
        \necount_RNO[1]_net_1 ));
    OR3C \timecount_RNO_5[18]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[18]_net_1 ), .Y(
        \OPENTIME_TEL_m[18] ));
    DFN1E0 \OPENTIME_TEL[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[0]_net_1 ));
    DFN1 \strippluse[1]  (.D(\strippluse_RNO[1]_net_1 ), .CLK(GLA), .Q(
        strippluse[1]));
    AOI1B \timecount_RNO_8[5]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[5]_net_1 ), .C(\CUTTIME180_TEL_m[5] ), .Y(
        \timecount_18_iv_3[5] ));
    OR2B \timecount_RNO_14[9]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[9]_net_1 ), .Y(\CUTTIME180_TEL_m[9] ));
    OR2 \CS_RNIPEHP[12]  (.A(N_1348), .B(N_1347), .Y(N_1393));
    NOR3C \timecount_RNO_2[10]  (.A(\OPENTIME_TEL_m[10] ), .B(
        \CUTTIME180_Tini_m[10] ), .C(\timecount_18_iv_3[10] ), .Y(
        \timecount_18_iv_7[10] ));
    NOR2 \CS_RNISJF6[1]  (.A(\CS[16]_net_1 ), .B(\CS[1]_net_1 ), .Y(
        N_1343));
    DFN1E1 \PLUSETIME180[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[13]_net_1 ));
    NOR2A \CS_RNO[5]  (.A(top_code_0_scale_rst), .B(N_1300), .Y(
        \CS_RNO_3[5] ));
    OR3C \timecount_RNO_7[4]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[4]_net_1 ), .Y(
        \ACQTIME_m[4] ));
    OR3C \timecount_RNO_7[10]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[10]_net_1 ), .Y(
        \OPENTIME_TEL_m[10] ));
    OR2 \CS_RNIH1N[14]  (.A(N_1344), .B(\CS[14]_net_1 ), .Y(N_1351));
    NOR2A \CS_RNO[14]  (.A(top_code_0_scale_rst), .B(N_1308), .Y(
        \CS_RNO[14]_net_1 ));
    OR3B CUTTIME180_Tini_265_e (.A(N_62), .B(
        un1_PLUSETIME9030_3_i_a2_0_net_1), .C(scalechoice[0]), .Y(
        N_1564_i));
    MX2 \strippluse_RNO_0[4]  (.A(\strippluse_6[4] ), .B(strippluse[4])
        , .S(un1_CS6_28), .Y(N_364));
    NOR2B intertodsp_RNO (.A(top_code_0_scale_rst), .B(N_508), .Y(
        intertodsp_RNO_0_net_1));
    OR2B \timecount_RNO_12[9]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[9]_net_1 ), .Y(\CUTTIME180_m[9] ));
    DFN1E0 \OPENTIME_TEL[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[10]_net_1 ));
    MX2C \strippluse_RNO_2[6]  (.A(\STRIPNUM90_NUM[6]_net_1 ), .B(
        \STRIPNUM180_NUM[6]_net_1 ), .S(\NS[8] ), .Y(N_242));
    AOI1B \timecount_RNO_9[1]  (.A(\S_DUMPTIME[1]_net_1 ), .B(
        N_1188_i_0), .C(\timecount_18_iv_10_2[1] ), .Y(
        \timecount_18_iv_10_6[1] ));
    NOR2B \strippluse_RNO[10]  (.A(top_code_0_scale_rst), .B(N_370), 
        .Y(\strippluse_RNO[10]_net_1 ));
    DFN1E1 \PLUSETIME90[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[15]_net_1 ));
    NOR2B \necount_RNO[3]  (.A(top_code_0_scale_rst), .B(N_514), .Y(
        \necount_RNO[3]_net_1 ));
    DFN1E1 \DUMPTIME[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[13]_net_1 ));
    MX2C \strippluse_RNO_2[3]  (.A(\STRIPNUM90_NUM[3]_net_1 ), .B(
        \STRIPNUM180_NUM[3]_net_1 ), .S(\NS[8] ), .Y(N_239));
    NOR2B \s_acqnum_1_RNO[10]  (.A(top_code_0_scale_rst), .B(N_358), 
        .Y(\s_acqnum_1_RNO[10]_net_1 ));
    OR3A intertodsp_RNO_2 (.A(N_1349), .B(N_1350), .C(\CS[16]_net_1 ), 
        .Y(N_1322));
    DFN1E1 \ACQTIME[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[5]_net_1 ));
    NOR2A \CS_RNO[7]  (.A(top_code_0_scale_rst), .B(N_1302), .Y(
        \CS_RNO_3[7] ));
    OR2B \timecount_RNO_6[7]  (.A(N_1185_i_0), .B(\DUMPTIME[7]_net_1 ), 
        .Y(\DUMPTIME_m[7] ));
    GND GND_i_0 (.Y(GND_0));
    NOR3 \CS_RNIG0OL[19]  (.A(timecount_12_sqmuxa), .B(N_1160_i_0), .C(
        N_1188_i_0), .Y(un1_timecount_5_sqmuxa_5));
    NOR2B s_acq_RNO (.A(top_code_0_scale_rst), .B(N_505), .Y(
        s_acq_RNO_0_net_1));
    DFN1E0 \OPENTIME[10]  (.D(scaledatain[10]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[10]_net_1 ));
    DFN1E1 \PLUSETIME90[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[4]_net_1 ));
    NOR2B \CS_RNI3LF1[12]  (.A(necount_LE_M_net_1), .B(\CS[12]_net_1 ), 
        .Y(timecount_11_sqmuxa_0));
    DFN1E1 \PLUSETIME90[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[10]_net_1 ));
    AOI1B \timecount_RNO_13[2]  (.A(\PLUSETIME180[2]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[2] ), .Y(\timecount_18_iv_1[2] )
        );
    NOR2A \CS_RNI3K7D[7]  (.A(\CS_i[0]_net_1 ), .B(\CS[7]_net_1 ), .Y(
        un1_CS6_39_i_a2_0));
    DFN1E0 \CUTTIME90[19]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1508), 
        .Q(\CUTTIME90[19]_net_1 ));
    DFN1E0 \OPENTIME[11]  (.D(scaledatain[11]), .CLK(GLA), .E(N_1436_i)
        , .Q(\OPENTIME[11]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[18]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[18]_net_1 ));
    OR2B \timecount_RNO_6[6]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[6]_net_1 ), .Y(\CUTTIME180_TEL_m[6] ));
    MX2 \s_acqnum_1_RNO_0[0]  (.A(\s_acqnum_7[0] ), .B(s_acqnum_1[0]), 
        .S(un1_CS6_28), .Y(N_348));
    DFN1E0 \CUTTIME180[3]  (.D(scaledatain[3]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[3]_net_1 ));
    NOR2A \CS_RNICUBC[10]  (.A(top_code_0_scale_rst), .B(N_1305), .Y(
        \CS_RNICUBC[10]_net_1 ));
    DFN1E0 \CUTTIME90[7]  (.D(scaledatain[7]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[7]_net_1 ));
    OR3C \timecount_RNO_12[5]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[5]_net_1 ), .Y(
        \ACQTIME_m[5] ));
    DFN1E1 \STRIPNUM90_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[2]_net_1 ));
    OR2B un1_PLUSETIME9030_i_a2_0 (.A(scalechoice[3]), .B(N_59), .Y(
        N_63));
    OR2B \timecount_RNO_12[7]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[7]_net_1 ), .Y(\CUTTIME180_m[7] ));
    DFN1E1 \NE_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[4]_net_1 ));
    DFN1E1 \STRIPNUM180_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[5]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[21]  (.D(scaledatain[5]), .CLK(GLA), .E(
        N_1596), .Q(\CUTTIME180_Tini[21]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[9]_net_1 ));
    DFN1E0 \CUTTIME180_Tini[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[0]_net_1 ));
    DFN1E1 \STRIPNUM90_NUM[6]  (.D(scaledatain[6]), .CLK(GLA), .E(
        STRIPNUM90_NUM_1_sqmuxa), .Q(\STRIPNUM90_NUM[6]_net_1 ));
    DFN1E1 \ACQ180_NUM[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[10]_net_1 ));
    DFN1E1 \M_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[2]_net_1 ));
    NOR2 \CS_RNILITK[14]  (.A(N_1392_i), .B(N_1351), .Y(N_1395));
    OR2B \timecount_RNO_9[13]  (.A(N_1185_i_0), .B(
        \DUMPTIME[13]_net_1 ), .Y(\DUMPTIME_m[13] ));
    OR3C \timecount_RNO[14]  (.A(\timecount_18_iv_4[14] ), .B(
        \timecount_18_iv_3[14] ), .C(\timecount_18_iv_8[14] ), .Y(
        \timecount_18[14] ));
    DFN1E1 \S_DUMPTIME[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[12]_net_1 ));
    DFN1 bb_ch (.D(bb_ch_RNO_net_1), .CLK(GLA), .Q(net_51));
    OR2B \timecount_RNO_3[19]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[19]_net_1 ), .Y(\CUTTIME180_TEL_m[19] ));
    MX2A \CS_RNO_0[1]  (.A(\CS[1]_net_1 ), .B(\CS_i[0]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1296));
    DFN1E1 \PLUSETIME180[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[4]_net_1 ));
    OR2B s_acq180_RNO_1 (.A(un1_CS6_0), .B(N_1278), .Y(un1_CS6));
    MX2C \strippluse_RNO_2[7]  (.A(\STRIPNUM90_NUM[7]_net_1 ), .B(
        \STRIPNUM180_NUM[7]_net_1 ), .S(\NS[8] ), .Y(N_243));
    DFN1 \strippluse[2]  (.D(\strippluse_RNO[2]_net_1 ), .CLK(GLA), .Q(
        strippluse[2]));
    DFN1E1 \ACQ180_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[2]_net_1 ));
    DFN1E1 \DUMPTIME[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[10]_net_1 ));
    OR2A sw_acq1_RNO (.A(top_code_0_scale_rst), .B(N_345), .Y(
        sw_acq1_RNO_0_net_1));
    NOR2B \strippluse_RNO[5]  (.A(top_code_0_scale_rst), .B(N_365), .Y(
        \strippluse_RNO[5]_net_1 ));
    NOR3C \timecount_RNO_4[4]  (.A(\OPENTIME_TEL_m[4] ), .B(
        \CUTTIME180_Tini_m[4] ), .C(\timecount_18_iv_3[4] ), .Y(
        \timecount_18_iv_7[4] ));
    XNOR2 M_pulse_RNO_8 (.A(\necount[2]_net_1 ), .B(\M_NUM[2]_net_1 ), 
        .Y(M_pulse8_2_i));
    DFN1E1 \ACQ180_NUM[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        ACQ180_NUM_1_sqmuxa), .Q(\ACQ180_NUM[8]_net_1 ));
    DFN1 dump_sustain_ctrl (.D(dump_sustain_ctrl_RNO_net_1), .CLK(GLA), 
        .Q(scalestate_0_dump_sustain_ctrl));
    AOI1B \timecount_RNO_1[16]  (.A(N_1162_i_0), .B(
        \CUTTIME90[16]_net_1 ), .C(\CUTTIME180_m[16] ), .Y(
        \timecount_18_0_iv_0[16] ));
    DFN1E1 \M_NUM[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[4]_net_1 ));
    OAI1 s_acq_RNO_1 (.A(N_1342), .B(un1_CS6_17_i_a3_0), .C(N_1278), 
        .Y(N_1259));
    OR3C \timecount_RNO_10[13]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[13]_net_1 ), .Y(
        \ACQTIME_m[13] ));
    OR3C \timecount_RNO[8]  (.A(\timecount_18_iv_4[8] ), .B(
        \timecount_18_iv_3[8] ), .C(\timecount_18_iv_8[8] ), .Y(
        \timecount_18[8] ));
    DFN1 \CS[5]  (.D(\CS_RNO_3[5] ), .CLK(GLA), .Q(\CS[5]_net_1 ));
    DFN1E1 \ACQTIME[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[14]_net_1 ));
    NOR2A \CS_RNO[15]  (.A(top_code_0_scale_rst), .B(N_1309), .Y(
        \CS_RNO[15]_net_1 ));
    XNOR2 fst_lst_pulse_RNO_6 (.A(\necount[5]_net_1 ), .B(
        \NE_NUM[5]_net_1 ), .Y(fst_lst_pulse8_5_i));
    OR3B \timecount_RNO_2[2]  (.A(top_code_0_scale_rst), .B(N_1328), 
        .C(\CS_RNITMND1[6]_net_1 ), .Y(\timecount_cnst_m[2] ));
    AOI1B \timecount_RNO_11[13]  (.A(\PLUSETIME180[13]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[13] ), .Y(
        \timecount_18_iv_1[13] ));
    OR2B \timecount_RNO_4[12]  (.A(N_1185_i_0), .B(
        \DUMPTIME[12]_net_1 ), .Y(\DUMPTIME_m[12] ));
    NOR2B \necount_RNO[2]  (.A(top_code_0_scale_rst), .B(N_513), .Y(
        \necount_RNO[2]_net_1 ));
    DFN1E1 \PLUSETIME180[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[11]_net_1 ));
    DFN1 s_acq (.D(s_acq_RNO_0_net_1), .CLK(GLA), .Q(
        scalestate_0_s_acq));
    MX2 \necount_RNO_0[9]  (.A(\necount1[9] ), .B(\necount[9]_net_1 ), 
        .S(N_1249), .Y(N_520));
    OR2A \necount_RNO[0]  (.A(top_code_0_scale_rst), .B(N_511), .Y(
        \necount_RNO[0]_net_1 ));
    NOR3C \timecount_RNO_4[9]  (.A(\OPENTIME_TEL_m[9] ), .B(
        \CUTTIME180_Tini_m[9] ), .C(timecount_18_iv_9_m1_e_3), .Y(
        timecount_18_iv_9_m1_e_7));
    OR2A fst_lst_pulse_RNI88CH (.A(N_1320), .B(fst_lst_pulse_net_1), 
        .Y(sw_acq1_1_sqmuxa));
    DFN1E0 \CUTTIME180_Tini[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[9]_net_1 ));
    OR2B \timecount_RNO_12[4]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[4]_net_1 ), .Y(\CUTTIME180_m[4] ));
    DFN1E1 \M_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[9]_net_1 ));
    OR2B \timecount_RNO_9[3]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[3]_net_1 ), .Y(\CUTTIME180_m[3] ));
    DFN1E1 \timecount[15]  (.D(\timecount_18[15] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[15]));
    OR3C \timecount_RNO_7[0]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[0]_net_1 ), .Y(
        \OPENTIME_TEL_m[0] ));
    OR3C CUTTIME180_197_e (.A(N_57), .B(N_62), .C(scalechoice[0]), .Y(
        N_1428));
    DFN1E1 \NE_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        NE_NUM_1_sqmuxa), .Q(\NE_NUM[0]_net_1 ));
    NOR3C M_pulse_RNO_3 (.A(M_pulse8_2_i), .B(M_pulse8_0_i), .C(
        M_pulse8_NE_1), .Y(M_pulse8_NE_6));
    NOR2B dump_sustain_ctrl_RNO (.A(top_code_0_scale_rst), .B(N_526), 
        .Y(dump_sustain_ctrl_RNO_net_1));
    DFN1E1 \M_NUM[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[5]_net_1 ));
    XNOR2 fst_lst_pulse_RNO_5 (.A(\necount[6]_net_1 ), .B(
        \NE_NUM[6]_net_1 ), .Y(fst_lst_pulse8_6_i));
    OR2B \timecount_RNO_6[9]  (.A(N_1185_i_0), .B(\DUMPTIME[9]_net_1 ), 
        .Y(\DUMPTIME_m[9] ));
    DFN1E0 \OPENTIME[4]  (.D(scaledatain[4]), .CLK(GLA), .E(N_1436_i), 
        .Q(\OPENTIME[4]_net_1 ));
    XNOR2 M_pulse_RNO_15 (.A(\necount[3]_net_1 ), .B(\M_NUM[3]_net_1 ), 
        .Y(M_pulse8_3_i));
    MX2C \CS_RNO_0[13]  (.A(\CS[13]_net_1 ), .B(\CS[12]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1307));
    AOI1B \timecount_RNO_2[19]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[19]_net_1 ), .C(\OPENTIME_TEL_m[19] ), .Y(
        \timecount_18_0_iv_2[19] ));
    DFN1E1 \timecount[21]  (.D(\timecount_18[21] ), .CLK(GLA), .E(
        un1_CS6_33), .Q(timecount[21]));
    DFN1E0 \CUTTIME180_TEL[18]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[18]_net_1 ));
    NOR2A \CS_RNO[10]  (.A(top_code_0_scale_rst), .B(N_1304), .Y(
        \CS_RNO[10]_net_1 ));
    NOR2A \CS_RNI360B[4]  (.A(top_code_0_scale_rst), .B(N_1346), .Y(
        N_1185_i_0));
    MX2 \s_acqnum_1_RNO_2[0]  (.A(\ACQ90_NUM[0]_net_1 ), .B(
        \ACQ180_NUM[0]_net_1 ), .S(\NS_0[8] ), .Y(N_264));
    DFN1E0 \CUTTIME180[6]  (.D(scaledatain[6]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[6]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[20]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1552), .Q(\CUTTIME180_TEL[20]_net_1 ));
    OR2 pn_out_RNO_1 (.A(top_code_0_pn_change), .B(\NS_0[8] ), .Y(
        un1_NS_2));
    AO1C \timecount_RNO[7]  (.A(\CS_RNITMND1[6]_net_1 ), .B(
        timecount_9_sqmuxa_m_0), .C(\timecount_18_iv_9[7] ), .Y(
        \timecount_18[7] ));
    OR2A \CS_RNI9KN6[15]  (.A(N_1346), .B(\CS[15]_net_1 ), .Y(N_1350));
    DFN1E0 \OPENTIME_TEL[19]  (.D(scaledatain[3]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[19]_net_1 ));
    DFN1 \necount[9]  (.D(\necount_RNO[9]_net_1 ), .CLK(GLA), .Q(
        \necount[9]_net_1 ));
    DFN1E0 \OPENTIME_TEL[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[12]_net_1 ));
    DFN1E1 \PLUSETIME90[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[12]_net_1 ));
    necount_cmp_1 necount_cmp_1 (.NE_NUM({\NE_NUM[11]_net_1 , 
        \NE_NUM[10]_net_1 , \NE_NUM[9]_net_1 , \NE_NUM[8]_net_1 , 
        \NE_NUM[7]_net_1 , \NE_NUM[6]_net_1 , \NE_NUM[5]_net_1 , 
        \NE_NUM[4]_net_1 , \NE_NUM[3]_net_1 , \NE_NUM[2]_net_1 , 
        \NE_NUM[1]_net_1 , \NE_NUM[0]_net_1 }), .necount({
        \necount[11]_net_1 , \necount[10]_net_1 , \necount[9]_net_1 , 
        \necount[8]_net_1 , \necount[7]_net_1 , \necount[6]_net_1 , 
        \necount[5]_net_1 , \necount[4]_net_1 , \necount[3]_net_1 , 
        \necount[2]_net_1 , \necount[1]_net_1 , \necount[0]_net_1 }), 
        .necount_LE_NE_1(necount_LE_NE_1));
    DFN1E1 \PLUSETIME180[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[14]_net_1 ));
    DFN1E1 \PLUSETIME90[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        PLUSETIME90_0_sqmuxa), .Q(\PLUSETIME90[14]_net_1 ));
    NOR2A ACQ90_NUM_1_sqmuxa_0_a2 (.A(ACQ90_NUM_1_sqmuxa_1), .B(N_63), 
        .Y(ACQ90_NUM_1_sqmuxa));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \strippluse_RNO_1[6]  (.A(N_242), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[6] ));
    OR2B \timecount_RNO_10[14]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[14]_net_1 ), .Y(\CUTTIME180_m[14] ));
    DFN1E1 \DUMPTIME[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[5]_net_1 ));
    AOI1B \timecount_RNO_0[17]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[17]_net_1 ), .C(\CUTTIME180_TEL_m[17] ), .Y(
        \timecount_18_0_iv_1[17] ));
    NOR3C fst_lst_pulse_RNO_2 (.A(fst_lst_pulse8_6_i), .B(
        fst_lst_pulse8_5_i), .C(fst_lst_pulse8_NE_3), .Y(
        fst_lst_pulse8_NE_7));
    MX2 \s_acqnum_1_RNO_0[9]  (.A(\s_acqnum_7[9] ), .B(s_acqnum_1[9]), 
        .S(un1_CS6_28), .Y(N_357));
    OR2A \CS_RNI6177[20]  (.A(N_1346), .B(timecount_18_iv_1_m3_e_1_1), 
        .Y(timecount_18_iv_1_m3_e_1));
    OR2B \timecount_RNO_11[14]  (.A(N_1162_i_0), .B(
        \CUTTIME90[14]_net_1 ), .Y(\CUTTIME90_m[14] ));
    OR3C \timecount_RNO_10[6]  (.A(\CS[14]_net_1 ), .B(
        top_code_0_scale_rst), .C(\ACQTIME[6]_net_1 ), .Y(
        \ACQTIME_m[6] ));
    OR3C \timecount_RNO[6]  (.A(\timecount_18_iv_8[6] ), .B(
        \timecount_18_iv_7[6] ), .C(\timecount_cnst_m[6] ), .Y(
        \timecount_18[6] ));
    MX2 \s_acqnum_1_RNO_0[8]  (.A(\s_acqnum_7[8] ), .B(s_acqnum_1[8]), 
        .S(un1_CS6_28), .Y(N_356));
    AOI1B \timecount_RNO_5[8]  (.A(N_1162_i_0), .B(
        \CUTTIME90[8]_net_1 ), .C(\CUTTIME180_m[8] ), .Y(
        \timecount_18_iv_2[8] ));
    XA1A M_pulse_RNO_13 (.A(\M_NUM[11]_net_1 ), .B(\necount[11]_net_1 )
        , .C(M_pulse8_10_i), .Y(M_pulse8_NE_5));
    DFN1E0 \CUTTIME180[0]  (.D(scaledatain[0]), .CLK(GLA), .E(N_1396_i)
        , .Q(\CUTTIME180[0]_net_1 ));
    DFN1E0 \CUTTIME180_TEL[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[2]_net_1 ));
    OR3C \timecount_RNO_14[6]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[6]_net_1 ), .Y(
        \OPENTIME_TEL_m[6] ));
    DFN1E1 \S_DUMPTIME[8]  (.D(scaledatain[8]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[8]_net_1 ));
    MX2 load_out_RNO_0 (.A(N_1393), .B(scalestate_0_load_out), .S(
        N_1253), .Y(N_501));
    DFN1E0 \OPENTIME_TEL[18]  (.D(scaledatain[2]), .CLK(GLA), .E(
        N_1640), .Q(\OPENTIME_TEL[18]_net_1 ));
    OR2 \CS_RNI07HC[3]  (.A(\CS[9]_net_1 ), .B(\CS[3]_net_1 ), .Y(
        N_1342));
    OAI1 reset_out_RNO_2 (.A(N_1392_i), .B(un1_CS6_39_i_a3_1), .C(
        timer_top_0_clk_en_scale), .Y(N_1245));
    DFN1E0 \CUTTIME90[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[10]_net_1 ));
    NOR3C necount_LE_M_RNIGRV5 (.A(\CS[15]_net_1 ), .B(
        necount_LE_M_net_1), .C(top_code_0_scale_rst), .Y(
        timecount_14_sqmuxa));
    NOR2B necount_LE_M_RNO (.A(top_code_0_scale_rst), .B(
        necount_LE_M_1), .Y(necount_LE_M_RNO_net_1));
    OR2B \timecount_RNO_9[8]  (.A(N_1185_i_0), .B(\DUMPTIME[8]_net_1 ), 
        .Y(\DUMPTIME_m[8] ));
    OR2B \timecount_RNO_15[2]  (.A(\PLUSETIME90[2]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[2] ));
    DFN1E1 \PLUSETIME180[5]  (.D(scaledatain[5]), .CLK(GLA), .E(
        PLUSETIME180_1_sqmuxa), .Q(\PLUSETIME180[5]_net_1 ));
    OR2A fst_lst_pulse_RNI242I (.A(\NS[8] ), .B(fst_lst_pulse_net_1), 
        .Y(s_acqnum_1_sqmuxa));
    DFN1E0 \CUTTIME90[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[12]_net_1 ));
    DFN1E1 \DUMPTIME[14]  (.D(scaledatain[14]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[14]_net_1 ));
    DFN1E0 \CUTTIME90[6]  (.D(scaledatain[6]), .CLK(GLA), .E(N_1476_i), 
        .Q(\CUTTIME90[6]_net_1 ));
    MX2C \CS_RNO_0[16]  (.A(\CS[16]_net_1 ), .B(\CS[15]_net_1 ), .S(
        timer_top_0_clk_en_scale_0), .Y(N_1310));
    NOR3A PLUSETIME90_0_sqmuxa_0_a2 (.A(N_59), .B(N_58), .C(
        scalechoice[0]), .Y(PLUSETIME90_0_sqmuxa));
    OR3C \timecount_RNO[18]  (.A(\timecount_18_0_iv_1[18] ), .B(
        \timecount_18_0_iv_0[18] ), .C(\timecount_18_0_iv_2[18] ), .Y(
        \timecount_18[18] ));
    NOR3 reset_out_RNO_1 (.A(un1_CS_32_0_a3_0), .B(\CS[16]_net_1 ), .C(
        \CS_0[11]_net_1 ), .Y(N_1323));
    DFN1E0 \OPENTIME_TEL[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[15]_net_1 ));
    DFN1 \strippluse[11]  (.D(\strippluse_RNO[11]_net_1 ), .CLK(GLA), 
        .Q(strippluse[11]));
    AOI1B \timecount_RNO_3[12]  (.A(N_1162_i_0), .B(
        \CUTTIME90[12]_net_1 ), .C(\CUTTIME180_m[12] ), .Y(
        \timecount_18_iv_2[12] ));
    NOR2B bb_ch_RNO (.A(top_code_0_scale_rst), .B(N_510), .Y(
        bb_ch_RNO_net_1));
    DFN1E1 \M_NUM[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        M_NUM_1_sqmuxa), .Q(\M_NUM[11]_net_1 ));
    OR2B dump_start_RNO_1 (.A(timer_top_0_clk_en_scale_0), .B(N_1319), 
        .Y(N_1251));
    DFN1E0 \CUTTIME180_Tini[1]  (.D(scaledatain[1]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[1]_net_1 ));
    OR3C fst_lst_pulse_RNI7OKG1 (.A(s_acqnum_1_sqmuxa), .B(N_1179), .C(
        N_1278), .Y(un1_CS6_28));
    AOI1B \timecount_RNO_8[7]  (.A(\PLUSETIME180[7]_net_1 ), .B(
        N_1156_i_0), .C(\PLUSETIME90_m[7] ), .Y(\timecount_18_iv_1[7] )
        );
    NOR3C un1_PLUSETIME9030_2_i_a2_0_0 (.A(top_code_0_scaleload), .B(
        scalechoice[4]), .C(scalechoice[1]), .Y(
        un1_PLUSETIME9030_3_i_a2_0_net_1));
    DFN1E1 \ACQECHO_NUM[0]  (.D(scaledatain[0]), .CLK(GLA), .E(
        ACQECHO_NUM_1_sqmuxa), .Q(\ACQECHO_NUM[0]_net_1 ));
    OR2B \timecount_RNO_8[15]  (.A(\PLUSETIME90[15]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[15] ));
    OR2B \timecount_RNO_5[1]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[1]_net_1 ), .Y(\CUTTIME180_Tini_m[1] ));
    XA1A M_pulse_RNO_10 (.A(\M_NUM[1]_net_1 ), .B(\necount[1]_net_1 ), 
        .C(M_pulse8_3_i), .Y(M_pulse8_NE_1));
    VCC VCC_i (.Y(VCC));
    OR2B \timecount_RNO_4[0]  (.A(N_1185_i_0), .B(\DUMPTIME[0]_net_1 ), 
        .Y(\DUMPTIME_m[0] ));
    OR3C \timecount_RNO[20]  (.A(\OPENTIME_TEL_m[20] ), .B(
        \CUTTIME180_Tini_m[20] ), .C(\timecount_18_0_iv_0[20] ), .Y(
        \timecount_18[20] ));
    AOI1B \timecount_RNO_1[11]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[11]_net_1 ), .C(\CUTTIME180_TEL_m[11] ), .Y(
        \timecount_18_iv_3[11] ));
    DFN1E1 \STRIPNUM180_NUM[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        STRIPNUM180_NUM_1_sqmuxa), .Q(\STRIPNUM180_NUM[9]_net_1 ));
    NOR3C \timecount_RNO_4[7]  (.A(\OPENTIME_TEL_m[7] ), .B(
        \CUTTIME180_Tini_m[7] ), .C(\timecount_18_iv_3[7] ), .Y(
        \timecount_18_iv_7[7] ));
    DFN1E0 \CUTTIME180_TEL[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[4]_net_1 ));
    AO1 \CS_RNIVM7D[7]  (.A(necount_LE_NE_net_1), .B(\CS[17]_net_1 ), 
        .C(\CS[7]_net_1 ), .Y(\NS[8] ));
    DFN1E0 \CUTTIME180[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[12]_net_1 ));
    AOI1B \timecount_RNO_0[15]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[15]_net_1 ), .C(\OPENTIME_TEL_m[15] ), .Y(
        \timecount_18_iv_4[15] ));
    XA1A fst_lst_pulse_RNO_10 (.A(\NE_NUM[1]_net_1 ), .B(
        \necount[1]_net_1 ), .C(fst_lst_pulse8_3_i), .Y(
        fst_lst_pulse8_NE_1));
    DFN1E0 \CUTTIME180_TEL[15]  (.D(scaledatain[15]), .CLK(GLA), .E(
        N_1520_i), .Q(\CUTTIME180_TEL[15]_net_1 ));
    DFN1E1 \S_DUMPTIME[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[2]_net_1 ));
    OR2B \timecount_RNO_3[21]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[21]_net_1 ), .Y(\CUTTIME180_TEL_m[21] ));
    DFN1E1 \ACQTIME[13]  (.D(scaledatain[13]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[13]_net_1 ));
    NOR2A \CS_RNO[6]  (.A(top_code_0_scale_rst), .B(N_1301), .Y(
        \CS_RNO_3[6] ));
    DFN1E0 \CUTTIME90[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        N_1476_i), .Q(\CUTTIME90[11]_net_1 ));
    MX2 \s_acqnum_1_RNO_0[2]  (.A(\s_acqnum_7[2] ), .B(s_acqnum_1[2]), 
        .S(un1_CS6_28), .Y(N_350));
    DFN1E1 \S_DUMPTIME[10]  (.D(scaledatain[10]), .CLK(GLA), .E(
        S_DUMPTIME_1_sqmuxa), .Q(\S_DUMPTIME[10]_net_1 ));
    NOR2 \strippluse_RNO_1[1]  (.A(N_237), .B(\CS[11]_net_1 ), .Y(
        \strippluse_6[1] ));
    DFN1E0 \CUTTIME180_Tini[12]  (.D(scaledatain[12]), .CLK(GLA), .E(
        N_1564_i), .Q(\CUTTIME180_Tini[12]_net_1 ));
    OR3C \timecount_RNO[10]  (.A(\timecount_18_iv_6[10] ), .B(
        \timecount_18_iv_5[10] ), .C(\timecount_18_iv_7[10] ), .Y(
        \timecount_18[10] ));
    OR2B \timecount_RNO_8[14]  (.A(\PLUSETIME90[14]_net_1 ), .B(
        N_1160_i_0), .Y(\PLUSETIME90_m[14] ));
    NOR3C \timecount_RNO_1[9]  (.A(timecount_18_iv_9_m1_e_6), .B(
        timecount_18_iv_9_m1_e_5), .C(timecount_18_iv_9_m1_e_7), .Y(
        timecount_18_iv_9_m1_e_9));
    NOR2A \CS_RNO[12]  (.A(top_code_0_scale_rst), .B(N_1306), .Y(
        \CS_RNO[12]_net_1 ));
    DFN1E1 \ACQTIME[9]  (.D(scaledatain[9]), .CLK(GLA), .E(
        ACQTIME_1_sqmuxa), .Q(\ACQTIME[9]_net_1 ));
    NOR3A un1_PLUSETIME9030_5_i_a2_0 (.A(top_code_0_scaleload), .B(
        scalechoice[4]), .C(scalechoice[1]), .Y(N_59));
    MX2 \s_acqnum_1_RNO_0[3]  (.A(\s_acqnum_7[3] ), .B(s_acqnum_1[3]), 
        .S(un1_CS6_28), .Y(N_351));
    NOR2B \necount_RNO[8]  (.A(top_code_0_scale_rst), .B(N_519), .Y(
        \necount_RNO[8]_net_1 ));
    XA1A M_pulse_RNO_7 (.A(\M_NUM[8]_net_1 ), .B(\necount[8]_net_1 ), 
        .C(M_pulse8_4_i), .Y(M_pulse8_NE_3));
    MX2 \s_acqnum_1_RNO_1[10]  (.A(N_274), .B(\ACQECHO_NUM[10]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[10] ));
    DFN1 \s_acqnum_1[6]  (.D(\s_acqnum_1_RNO[6]_net_1 ), .CLK(GLA), .Q(
        s_acqnum_1[6]));
    OR3C \timecount_RNO[12]  (.A(\timecount_18_iv_6[12] ), .B(
        \timecount_18_iv_5[12] ), .C(\timecount_18_iv_7[12] ), .Y(
        \timecount_18[12] ));
    MX2 \strippluse_RNO_0[0]  (.A(\strippluse_6[0] ), .B(strippluse[0])
        , .S(un1_CS6_28), .Y(N_360));
    NOR3C \timecount_RNO_5[5]  (.A(\DUMPTIME_m[5] ), .B(\ACQTIME_m[5] )
        , .C(\timecount_18_iv_1[5] ), .Y(\timecount_18_iv_5[5] ));
    OR2B \timecount_RNO_1[21]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[21]_net_1 ), .Y(\CUTTIME180_Tini_m[21] ));
    OR3 reset_out_RNO_4 (.A(\CS_0[11]_net_1 ), .B(\CS[6]_net_1 ), .C(
        N_1348), .Y(un1_CS6_39_i_a3_1));
    XNOR2 fst_lst_pulse_RNO_14 (.A(\necount[4]_net_1 ), .B(
        \NE_NUM[4]_net_1 ), .Y(fst_lst_pulse8_4_i));
    MX2C \CS_RNO_0[12]  (.A(\CS[12]_net_1 ), .B(\CS[11]_net_1 ), .S(
        timer_top_0_clk_en_scale), .Y(N_1306));
    DFN1E1 \ACQ90_NUM[2]  (.D(scaledatain[2]), .CLK(GLA), .E(
        ACQ90_NUM_1_sqmuxa), .Q(\ACQ90_NUM[2]_net_1 ));
    OR3C \timecount_RNO_0[21]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[21]_net_1 ), .Y(
        \OPENTIME_TEL_m[21] ));
    NOR2 \strippluse_RNO_1[10]  (.A(N_246), .B(\CS_0[11]_net_1 ), .Y(
        \strippluse_6[10] ));
    NOR3C \timecount_RNO_1[2]  (.A(\OPENTIME_TEL_m[2] ), .B(
        \CUTTIME180_Tini_m[2] ), .C(\timecount_18_iv_3[2] ), .Y(
        \timecount_18_iv_7[2] ));
    DFN1 \CS[1]  (.D(\CS_RNO_3[1] ), .CLK(GLA), .Q(\CS[1]_net_1 ));
    AOI1B \timecount_RNO_0[14]  (.A(timecount_15_sqmuxa), .B(
        \CUTTIME180_Tini[14]_net_1 ), .C(\OPENTIME_TEL_m[14] ), .Y(
        \timecount_18_iv_4[14] ));
    MX2 \s_acqnum_1_RNO_1[0]  (.A(N_264), .B(\ACQECHO_NUM[0]_net_1 ), 
        .S(\CS_0[11]_net_1 ), .Y(\s_acqnum_7[0] ));
    DFN1E1 \DUMPTIME[7]  (.D(scaledatain[7]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa), .Q(\DUMPTIME[7]_net_1 ));
    NOR3C \timecount_RNO_3[4]  (.A(\DUMPTIME_m[4] ), .B(\ACQTIME_m[4] )
        , .C(\timecount_18_iv_1[4] ), .Y(\timecount_18_iv_5[4] ));
    OR2B \timecount_RNO_4[13]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[13]_net_1 ), .Y(\CUTTIME180_TEL_m[13] ));
    NOR3C \timecount_RNO_2[12]  (.A(\OPENTIME_TEL_m[12] ), .B(
        \CUTTIME180_Tini_m[12] ), .C(\timecount_18_iv_3[12] ), .Y(
        \timecount_18_iv_7[12] ));
    DFN1E0 \OPENTIME_TEL[4]  (.D(scaledatain[4]), .CLK(GLA), .E(
        N_1608_i), .Q(\OPENTIME_TEL[4]_net_1 ));
    AOI1B \timecount_RNO_9[0]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[0]_net_1 ), .C(\OPENTIME_m[0] ), .Y(
        \timecount_18_iv_3[0] ));
    OR2B \timecount_RNO_10[1]  (.A(timecount_14_sqmuxa), .B(
        \CUTTIME180_TEL[1]_net_1 ), .Y(\CUTTIME180_TEL_m[1] ));
    AOI1B \timecount_RNO_6[15]  (.A(N_1185_i_0), .B(
        \DUMPTIME[15]_net_1 ), .C(\ACQTIME_m[15] ), .Y(
        \timecount_18_iv_0[15] ));
    NOR2A \CS_RNO[1]  (.A(top_code_0_scale_rst), .B(N_1296), .Y(
        \CS_RNO_3[1] ));
    OR3C \timecount_RNO_7[12]  (.A(timecount_11_sqmuxa_0), .B(
        top_code_0_scale_rst), .C(\OPENTIME_TEL[12]_net_1 ), .Y(
        \OPENTIME_TEL_m[12] ));
    DFN1E0 \CUTTIME180[11]  (.D(scaledatain[11]), .CLK(GLA), .E(
        N_1396_i), .Q(\CUTTIME180[11]_net_1 ));
    NOR3C \timecount_RNO_1[10]  (.A(\DUMPTIME_m[10] ), .B(
        \ACQTIME_m[10] ), .C(\timecount_18_iv_1[10] ), .Y(
        \timecount_18_iv_5[10] ));
    OR2B \timecount_RNO_14[1]  (.A(timecount_16_sqmuxa), .B(
        \CUTTIME180[1]_net_1 ), .Y(\CUTTIME180_m[1] ));
    AOI1B \timecount_RNO_11[4]  (.A(timecount_12_sqmuxa), .B(
        \OPENTIME[4]_net_1 ), .C(\CUTTIME180_TEL_m[4] ), .Y(
        \timecount_18_iv_3[4] ));
    MX2 \s_acqnum_1_RNO_2[9]  (.A(\ACQ90_NUM[9]_net_1 ), .B(
        \ACQ180_NUM[9]_net_1 ), .S(\NS[8] ), .Y(N_273));
    
endmodule


module topctrlchange(
       change,
       GLA,
       plusestate_0_sw_acq1,
       scalestate_0_sw_acq1,
       plusestate_0_state_over_n,
       scalestate_0_tetw_pluse,
       nsctrl_choice_0_intertodsp,
       scalestate_0_sw_acq2,
       nsctrl_choice_0_sw_acq2,
       plusestate_0_soft_d,
       scalestate_0_soft_d,
       nsctrl_choice_0_soft_d,
       scalestate_0_rt_sw,
       nsctrl_choice_0_rt_sw,
       net_27,
       rt_sw_net_1,
       soft_dump_net_1,
       sw_acq1_c,
       sw_acq2_c,
       un1_change_2,
       interupt_c
    );
input  [1:0] change;
input  GLA;
input  plusestate_0_sw_acq1;
input  scalestate_0_sw_acq1;
input  plusestate_0_state_over_n;
input  scalestate_0_tetw_pluse;
input  nsctrl_choice_0_intertodsp;
input  scalestate_0_sw_acq2;
input  nsctrl_choice_0_sw_acq2;
input  plusestate_0_soft_d;
input  scalestate_0_soft_d;
input  nsctrl_choice_0_soft_d;
input  scalestate_0_rt_sw;
input  nsctrl_choice_0_rt_sw;
input  net_27;
output rt_sw_net_1;
output soft_dump_net_1;
output sw_acq1_c;
output sw_acq2_c;
input  un1_change_2;
output interupt_c;

    wire \un1_interin1[0] , interin3_m, interin2_m, interin1_m, 
        soft_dump_6, s_dumpin3_m, s_dumpin2_m, s_dumpin1_m, N_8, N_9, 
        sw_acq2_6_iv, N_10, sw_acq1_6_iv, N_11, N_12, rt_sw_6, 
        rt_sw_RNO_3, soft_dump_RNO_0_net_1, interupt_RNO_net_1, 
        sw_acq1_RNO_net_1, sw_acq2_RNO_2_net_1, rt_swin1_m, 
        sw_acq2in1_i_m, sw_acq1in2_i_m, GND, VCC, GND_0, VCC_0;
    
    OR3A soft_dump_RNO_4 (.A(nsctrl_choice_0_soft_d), .B(change[0]), 
        .C(change[1]), .Y(s_dumpin1_m));
    OA1C sw_acq1_RNO_1 (.A(change[1]), .B(plusestate_0_sw_acq1), .C(
        sw_acq1in2_i_m), .Y(sw_acq1_6_iv));
    NOR2B rt_sw_RNO (.A(N_12), .B(net_27), .Y(rt_sw_RNO_3));
    NOR2B interupt_RNO (.A(N_8), .B(net_27), .Y(interupt_RNO_net_1));
    MX2 sw_acq2_RNO_0 (.A(sw_acq2_c), .B(sw_acq2_6_iv), .S(
        un1_change_2), .Y(N_9));
    AO1B rt_sw_RNO_1 (.A(change[0]), .B(scalestate_0_rt_sw), .C(
        rt_swin1_m), .Y(rt_sw_6));
    NOR2B interupt_RNO_2 (.A(change[1]), .B(plusestate_0_state_over_n), 
        .Y(interin3_m));
    DFN1 sw_acq1 (.D(sw_acq1_RNO_net_1), .CLK(GLA), .Q(sw_acq1_c));
    VCC VCC_i (.Y(VCC));
    OA1C sw_acq2_RNO_1 (.A(change[0]), .B(scalestate_0_sw_acq2), .C(
        sw_acq2in1_i_m), .Y(sw_acq2_6_iv));
    MX2 sw_acq1_RNO_0 (.A(sw_acq1_c), .B(sw_acq1_6_iv), .S(
        un1_change_2), .Y(N_10));
    OR2B soft_dump_RNO_2 (.A(change[1]), .B(plusestate_0_soft_d), .Y(
        s_dumpin3_m));
    DFN1 rt_sw (.D(rt_sw_RNO_3), .CLK(GLA), .Q(rt_sw_net_1));
    DFN1 soft_dump (.D(soft_dump_RNO_0_net_1), .CLK(GLA), .Q(
        soft_dump_net_1));
    OR2A sw_acq1_RNO (.A(net_27), .B(N_10), .Y(sw_acq1_RNO_net_1));
    OR3C soft_dump_RNO_1 (.A(s_dumpin3_m), .B(s_dumpin2_m), .C(
        s_dumpin1_m), .Y(soft_dump_6));
    NOR2B interupt_RNO_3 (.A(change[0]), .B(scalestate_0_tetw_pluse), 
        .Y(interin2_m));
    NOR3 sw_acq2_RNO_2 (.A(change[0]), .B(change[1]), .C(
        nsctrl_choice_0_sw_acq2), .Y(sw_acq2in1_i_m));
    OR3A rt_sw_RNO_2 (.A(nsctrl_choice_0_rt_sw), .B(change[0]), .C(
        change[1]), .Y(rt_swin1_m));
    GND GND_i (.Y(GND));
    NOR3A interupt_RNO_4 (.A(nsctrl_choice_0_intertodsp), .B(change[0])
        , .C(change[1]), .Y(interin1_m));
    DFN1 sw_acq2 (.D(sw_acq2_RNO_2_net_1), .CLK(GLA), .Q(sw_acq2_c));
    OR2B soft_dump_RNO_3 (.A(change[0]), .B(scalestate_0_soft_d), .Y(
        s_dumpin2_m));
    NOR2B soft_dump_RNO (.A(N_11), .B(net_27), .Y(
        soft_dump_RNO_0_net_1));
    OR2A sw_acq2_RNO (.A(net_27), .B(N_9), .Y(sw_acq2_RNO_2_net_1));
    MX2 interupt_RNO_0 (.A(interupt_c), .B(\un1_interin1[0] ), .S(
        un1_change_2), .Y(N_8));
    MX2 soft_dump_RNO_0 (.A(soft_dump_net_1), .B(soft_dump_6), .S(
        un1_change_2), .Y(N_11));
    DFN1 interupt (.D(interupt_RNO_net_1), .CLK(GLA), .Q(interupt_c));
    MX2 rt_sw_RNO_0 (.A(rt_sw_net_1), .B(rt_sw_6), .S(un1_change_2), 
        .Y(N_12));
    NOR2A sw_acq1_RNO_2 (.A(change[0]), .B(scalestate_0_sw_acq1), .Y(
        sw_acq1in2_i_m));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR3 interupt_RNO_1 (.A(interin3_m), .B(interin2_m), .C(interin1_m)
        , .Y(\un1_interin1[0] ));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module xwe_xzcs2_syn(
       GLA,
       GPMI_0_code_en,
       xwe_c,
       net_27,
       zcs2_c
    );
input  GLA;
output GPMI_0_code_en;
input  xwe_c;
input  net_27;
input  zcs2_c;

    wire code_en_0_0, xwe_reg2_net_1, code_en_RNO_net_1, 
        xwe_reg1_net_1, xwe_reg2_RNO_net_1, xwe_reg1_RNO_net_1, GND, 
        VCC, GND_0, VCC_0;
    
    NOR3B code_en_RNO (.A(xwe_reg1_net_1), .B(net_27), .C(code_en_0_0), 
        .Y(code_en_RNO_net_1));
    OR2 code_en_RNO_0 (.A(zcs2_c), .B(xwe_reg2_net_1), .Y(code_en_0_0));
    DFN1 code_en (.D(code_en_RNO_net_1), .CLK(GLA), .Q(GPMI_0_code_en));
    DFN1 xwe_reg2 (.D(xwe_reg2_RNO_net_1), .CLK(GLA), .Q(
        xwe_reg2_net_1));
    NOR2B xwe_reg2_RNO (.A(net_27), .B(xwe_reg1_net_1), .Y(
        xwe_reg2_RNO_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    VCC VCC_i (.Y(VCC));
    NOR2B xwe_reg1_RNO (.A(xwe_c), .B(net_27), .Y(xwe_reg1_RNO_net_1));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    DFN1 xwe_reg1 (.D(xwe_reg1_RNO_net_1), .CLK(GLA), .Q(
        xwe_reg1_net_1));
    
endmodule


module tri_state(
       zcs2_c,
       tri_ctrl_c,
       xd_1
    );
input  zcs2_c;
input  tri_ctrl_c;
output xd_1;

    wire GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    NOR2A xd_1_inst_1 (.A(tri_ctrl_c), .B(zcs2_c), .Y(xd_1));
    GND GND_i (.Y(GND));
    
endmodule


module rst_n_module(
       rst_n_module_VCC,
       INV_0_Y,
       GLA,
       net_27
    );
input  rst_n_module_VCC;
input  INV_0_Y;
input  GLA;
output net_27;

    wire rst_nr2_net_1, rst_nr1_net_1, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1C0 rst_nr1 (.D(rst_n_module_VCC), .CLK(GLA), .CLR(INV_0_Y), .Q(
        rst_nr1_net_1));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    CLKINT rst_nr2_RNIODQ1 (.A(rst_nr2_net_1), .Y(net_27));
    DFN1C0 rst_nr2 (.D(rst_nr1_net_1), .CLK(GLA), .CLR(INV_0_Y), .Q(
        rst_nr2_net_1));
    GND GND_i (.Y(GND));
    
endmodule


module GPMI(
       GPMI_VCC,
       xd_1,
       tri_ctrl_c,
       zcs2_c,
       net_27,
       xwe_c,
       GPMI_0_code_en,
       GLA,
       gpio_c
    );
input  GPMI_VCC;
output xd_1;
input  tri_ctrl_c;
input  zcs2_c;
output net_27;
input  xwe_c;
output GPMI_0_code_en;
input  GLA;
input  gpio_c;

    wire INV_0_Y, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    INV INV_0 (.A(gpio_c), .Y(INV_0_Y));
    xwe_xzcs2_syn xwe_xzcs2_syn_0 (.GLA(GLA), .GPMI_0_code_en(
        GPMI_0_code_en), .xwe_c(xwe_c), .net_27(net_27), .zcs2_c(
        zcs2_c));
    VCC VCC_i (.Y(VCC));
    tri_state tri_state_0 (.zcs2_c(zcs2_c), .tri_ctrl_c(tri_ctrl_c), 
        .xd_1(xd_1));
    rst_n_module rst_n_module_0 (.rst_n_module_VCC(GPMI_VCC), .INV_0_Y(
        INV_0_Y), .GLA(GLA), .net_27(net_27));
    GND GND_i (.Y(GND));
    
endmodule


module plusestate(
       timecount_1_1,
       plusedata,
       GLA,
       plusestate_0_off_test,
       plusestate_0_sw_acq1,
       plusestate_0_pluse_acq,
       plusestate_0_dds_config,
       plusestate_0_state_over_n,
       top_code_0_pluse_rst,
       top_code_0_pluse_lc,
       top_code_0_pluseload,
       plusestate_0_tetw_pluse,
       timer_top_0_clk_en_pluse,
       plusestate_0_soft_d,
       top_code_0_pluse_rst_0
    );
output [15:0] timecount_1_1;
input  [15:0] plusedata;
input  GLA;
output plusestate_0_off_test;
output plusestate_0_sw_acq1;
output plusestate_0_pluse_acq;
output plusestate_0_dds_config;
output plusestate_0_state_over_n;
input  top_code_0_pluse_rst;
input  top_code_0_pluse_lc;
input  top_code_0_pluseload;
output plusestate_0_tetw_pluse;
input  timer_top_0_clk_en_pluse;
output plusestate_0_soft_d;
input  top_code_0_pluse_rst_0;

    wire \timecount_5_i_1[7] , \PLUSETIME[7]_net_1 , N_153, 
        \timecount_5_i_0[7] , \DUMPTIME[7]_net_1 , \CS[5]_net_1 , 
        \timecount_5_i_1[2] , \PLUSETIME[2]_net_1 , 
        \timecount_5_i_0[2] , \DUMPTIME[2]_net_1 , 
        \timecount_5_i_1[4] , \PLUSETIME[4]_net_1 , 
        \timecount_5_i_0[4] , \DUMPTIME[4]_net_1 , 
        \timecount_5_i_1[5] , \PLUSETIME[5]_net_1 , 
        \timecount_5_i_0[5] , \DUMPTIME[5]_net_1 , 
        \timecount_5_i_0[6] , \DUMPTIME[6]_net_1 , 
        \timecount_5_i_0[8] , \DUMPTIME[8]_net_1 , 
        \timecount_5_i_0[1] , \DUMPTIME[1]_net_1 , 
        \timecount_5_i_0[3] , \DUMPTIME[3]_net_1 , 
        \timecount_5_1_0[0] , \DUMPTIME[0]_net_1 , N_19, N_140, N_155, 
        N_15, N_135, N_156, N_13, \CS[4]_net_1 , N_11, \CS[3]_net_1 , 
        N_7, \timecount_5[0] , \PLUSETIME[0]_net_1 , N_351, N_354, 
        N_92, N_116, \CS_i[0]_net_1 , N_152, N_5, N_115, N_350, 
        \CS[8]_net_1 , N_9, N_120, N_122, N_17, N_125, 
        \PLUSETIME[6]_net_1 , \PLUSETIME[8]_net_1 , \CS[9]_net_1 , 
        N_23, N_97, N_71, N_25, N_98, N_27, N_99, N_31, N_101, N_33, 
        N_102, \CS_RNO[1]_net_1 , N_103, \CS_RNO[2]_net_1 , N_104, 
        \CS_RNO[5]_net_1 , N_107, \CS_RNO[6]_net_1 , N_108, 
        \CS_i_RNO[0]_net_1 , N_61, N_65, N_91, \CS[2]_net_1 , 
        \CS[1]_net_1 , \PLUSETIME[10]_net_1 , \DUMPTIME[10]_net_1 , 
        \PLUSETIME[11]_net_1 , \DUMPTIME[11]_net_1 , 
        \PLUSETIME[12]_net_1 , \DUMPTIME[12]_net_1 , 
        \PLUSETIME[14]_net_1 , \DUMPTIME[14]_net_1 , 
        \PLUSETIME[15]_net_1 , \DUMPTIME[15]_net_1 , \CS[6]_net_1 , 
        DUMPTIME_1_sqmuxa_net_1, DUMPTIME_0_sqmuxa_net_1, 
        \PLUSETIME[1]_net_1 , \CS_RNO[7]_net_1 , \CS[7]_net_1 , 
        un1_sw_acq1_2_sqmuxa, N_109, N_106, N_105, 
        state_over_n_RNO_net_1, N_63, N_126, N_57, N_146, 
        \CS_RNO[8]_net_1 , \CS_RNO[4]_net_1 , \CS_RNO[3]_net_1 , N_357, 
        N_151, N_124, \PLUSETIME[3]_net_1 , N_110, N_100, 
        \PLUSETIME[13]_net_1 , \DUMPTIME[13]_net_1 , N_96, 
        \PLUSETIME[9]_net_1 , \DUMPTIME[9]_net_1 , N_59, N_145, 
        \CS_RNO[9]_net_1 , N_29, N_21, GND, VCC, GND_0, VCC_0;
    
    OA1B \timecount_1_RNO_0[3]  (.A(\CS[8]_net_1 ), .B(N_91), .C(N_152)
        , .Y(N_120));
    MX2C \timecount_1_RNO_0[12]  (.A(\PLUSETIME[12]_net_1 ), .B(
        \DUMPTIME[12]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_99));
    NOR2 \timecount_1_RNO[10]  (.A(N_97), .B(N_71), .Y(N_23));
    DFN1E1 \timecount_1[0]  (.D(\timecount_5[0] ), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[0]));
    DFN1E1 \PLUSETIME[12]  (.D(plusedata[12]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[12]_net_1 ));
    DFN1E1 \timecount_1[1]  (.D(N_5), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[1]));
    OR2A \CS_RNIKNR7[9]  (.A(\CS[9]_net_1 ), .B(\CS[5]_net_1 ), .Y(
        N_153));
    DFN1E1 \PLUSETIME[11]  (.D(plusedata[11]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[11]_net_1 ));
    DFN1E1 \PLUSETIME[9]  (.D(plusedata[9]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[9]_net_1 ));
    NOR2A \CS_RNO[4]  (.A(top_code_0_pluse_rst), .B(N_106), .Y(
        \CS_RNO[4]_net_1 ));
    OA1B \timecount_1_RNO[5]  (.A(\CS[4]_net_1 ), .B(N_156), .C(
        \timecount_5_i_1[5] ), .Y(N_13));
    NOR2A \CS_RNO[9]  (.A(top_code_0_pluse_rst), .B(N_110), .Y(
        \CS_RNO[9]_net_1 ));
    DFN1E1 \DUMPTIME[12]  (.D(plusedata[12]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[12]_net_1 ));
    NOR2A DUMPTIME_0_sqmuxa (.A(top_code_0_pluseload), .B(
        top_code_0_pluse_lc), .Y(DUMPTIME_0_sqmuxa_net_1));
    OA1B \timecount_1_RNO[7]  (.A(\CS[4]_net_1 ), .B(N_155), .C(
        \timecount_5_i_1[7] ), .Y(N_17));
    DFN1 \CS[4]  (.D(\CS_RNO[4]_net_1 ), .CLK(GLA), .Q(\CS[4]_net_1 ));
    OA1A \timecount_1_RNO_1[8]  (.A(\CS[5]_net_1 ), .B(
        \DUMPTIME[8]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[8] ));
    DFN1E1 \DUMPTIME[2]  (.D(plusedata[2]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[2]_net_1 ));
    MX2C \CS_RNO_0[4]  (.A(\CS[4]_net_1 ), .B(\CS[3]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_106));
    DFN1E1 \timecount_1[13]  (.D(N_29), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[13]));
    DFN1E1 \timecount_1[10]  (.D(N_23), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[10]));
    NOR3C \timecount_1_RNO[6]  (.A(N_135), .B(\timecount_5_i_0[6] ), 
        .C(N_156), .Y(N_15));
    MX2C \timecount_1_RNO_0[9]  (.A(\PLUSETIME[9]_net_1 ), .B(
        \DUMPTIME[9]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_96));
    DFN1E1 \PLUSETIME[14]  (.D(plusedata[14]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[14]_net_1 ));
    DFN1E1 \timecount_1[2]  (.D(N_7), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[2]));
    DFN1E1 \PLUSETIME[5]  (.D(plusedata[5]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[5]_net_1 ));
    MX2 soft_d_RNO_0 (.A(N_354), .B(plusestate_0_soft_d), .S(N_351), 
        .Y(N_125));
    DFN1E1 \DUMPTIME[4]  (.D(plusedata[4]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[4]_net_1 ));
    DFN1 \CS[3]  (.D(\CS_RNO[3]_net_1 ), .CLK(GLA), .Q(\CS[3]_net_1 ));
    MX2A sw_acq1_RNO_0 (.A(N_354), .B(plusestate_0_sw_acq1), .S(N_350), 
        .Y(N_124));
    DFN1E1 \DUMPTIME[1]  (.D(plusedata[1]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[1]_net_1 ));
    DFN1E1 \timecount_1[12]  (.D(N_27), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[12]));
    DFN1E1 \DUMPTIME[7]  (.D(plusedata[7]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[7]_net_1 ));
    DFN1E1 \DUMPTIME[9]  (.D(plusedata[9]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[9]_net_1 ));
    NOR2A \CS_RNO[5]  (.A(top_code_0_pluse_rst_0), .B(N_107), .Y(
        \CS_RNO[5]_net_1 ));
    MX2C \CS_RNO_0[5]  (.A(\CS[5]_net_1 ), .B(\CS[9]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_107));
    AO1D \timecount_1_RNO_0[5]  (.A(\PLUSETIME[5]_net_1 ), .B(N_153), 
        .C(\timecount_5_i_0[5] ), .Y(\timecount_5_i_1[5] ));
    DFN1E1 \PLUSETIME[15]  (.D(plusedata[15]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[15]_net_1 ));
    MX2A \CS_RNO_0[1]  (.A(\CS[1]_net_1 ), .B(\CS_i[0]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_103));
    DFN1E1 \timecount_1[8]  (.D(N_19), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[8]));
    NOR2B pluse_acq_RNO (.A(top_code_0_pluse_rst), .B(N_126), .Y(N_63));
    MX2C \timecount_1_RNO_0[10]  (.A(\PLUSETIME[10]_net_1 ), .B(
        \DUMPTIME[10]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_97));
    DFN1E1 \PLUSETIME[8]  (.D(plusedata[8]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[8]_net_1 ));
    OR2A sw_acq1_RNO (.A(top_code_0_pluse_rst), .B(N_124), .Y(N_151));
    DFN1E1 \DUMPTIME[8]  (.D(plusedata[8]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[8]_net_1 ));
    DFN1 \CS[1]  (.D(\CS_RNO[1]_net_1 ), .CLK(GLA), .Q(\CS[1]_net_1 ));
    GND GND_i (.Y(GND));
    AO1C \timecount_1_RNO_1[5]  (.A(\DUMPTIME[5]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[5] ));
    AO1C \timecount_1_RNO_1[2]  (.A(\DUMPTIME[2]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[2] ));
    DFN1E1 \PLUSETIME[10]  (.D(plusedata[10]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[10]_net_1 ));
    DFN1E1 \DUMPTIME[6]  (.D(plusedata[6]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[6]_net_1 ));
    OA1 \CS_i_RNO[0]  (.A(\CS_i[0]_net_1 ), .B(
        timer_top_0_clk_en_pluse), .C(top_code_0_pluse_rst_0), .Y(
        \CS_i_RNO[0]_net_1 ));
    DFN1 \CS_i[0]  (.D(\CS_i_RNO[0]_net_1 ), .CLK(GLA), .Q(
        \CS_i[0]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    AO1D \timecount_1_RNO_0[4]  (.A(\PLUSETIME[4]_net_1 ), .B(N_153), 
        .C(\timecount_5_i_0[4] ), .Y(\timecount_5_i_1[4] ));
    AO1D \timecount_1_RNO_0[2]  (.A(\PLUSETIME[2]_net_1 ), .B(N_153), 
        .C(\timecount_5_i_0[2] ), .Y(\timecount_5_i_1[2] ));
    OA1B \CS_RNO[7]  (.A(\CS[7]_net_1 ), .B(timer_top_0_clk_en_pluse), 
        .C(un1_sw_acq1_2_sqmuxa), .Y(\CS_RNO[7]_net_1 ));
    OR2 pluse_acq_RNO_1 (.A(N_92), .B(\CS[9]_net_1 ), .Y(N_357));
    OA1B \timecount_1_RNO[4]  (.A(\CS[3]_net_1 ), .B(N_155), .C(
        \timecount_5_i_1[4] ), .Y(N_11));
    NOR2B off_test_RNO (.A(top_code_0_pluse_rst), .B(N_145), .Y(N_59));
    DFN1E1 \timecount_1[11]  (.D(N_25), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[11]));
    NOR2B soft_d_RNO (.A(top_code_0_pluse_rst_0), .B(N_125), .Y(N_65));
    DFN1E1 \PLUSETIME[3]  (.D(plusedata[3]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[3]_net_1 ));
    DFN1E1 \timecount_1[5]  (.D(N_13), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[5]));
    NOR2A \CS_RNO[3]  (.A(top_code_0_pluse_rst), .B(N_105), .Y(
        \CS_RNO[3]_net_1 ));
    DFN1E1 \timecount_1[14]  (.D(N_31), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[14]));
    DFN1E1 \PLUSETIME[4]  (.D(plusedata[4]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[4]_net_1 ));
    DFN1 soft_d (.D(N_65), .CLK(GLA), .Q(plusestate_0_soft_d));
    MX2C \CS_RNO_0[6]  (.A(\CS[6]_net_1 ), .B(\CS[5]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_108));
    AO1C \timecount_1_RNO_1[4]  (.A(\DUMPTIME[4]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[4] ));
    DFN1 state_over_n (.D(state_over_n_RNO_net_1), .CLK(GLA), .Q(
        plusestate_0_state_over_n));
    NOR2A \CS_RNO[1]  (.A(top_code_0_pluse_rst_0), .B(N_103), .Y(
        \CS_RNO[1]_net_1 ));
    NOR3 \timecount_1_RNO[3]  (.A(N_120), .B(\timecount_5_i_0[3] ), .C(
        N_122), .Y(N_9));
    DFN1 \CS[9]  (.D(\CS_RNO[9]_net_1 ), .CLK(GLA), .Q(\CS[9]_net_1 ));
    VCC VCC_i (.Y(VCC));
    DFN1E1 \timecount_1[7]  (.D(N_17), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[7]));
    MX2C \CS_RNO_0[2]  (.A(\CS[2]_net_1 ), .B(\CS[1]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_104));
    NOR2 \timecount_1_RNO[12]  (.A(N_99), .B(N_71), .Y(N_27));
    DFN1E1 \timecount_1[15]  (.D(N_33), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[15]));
    OR2B \CS_RNI1K4E[9]  (.A(top_code_0_pluse_rst), .B(N_152), .Y(N_71)
        );
    NOR3A \timecount_1_RNO_0[1]  (.A(\CS_i[0]_net_1 ), .B(
        \CS[3]_net_1 ), .C(N_152), .Y(N_116));
    DFN1E1 \DUMPTIME[10]  (.D(plusedata[10]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[10]_net_1 ));
    AO1A dds_config_RNO_0 (.A(\CS[9]_net_1 ), .B(
        plusestate_0_dds_config), .C(N_92), .Y(N_146));
    AO1 pluse_acq_RNO_0 (.A(plusestate_0_pluse_acq), .B(N_354), .C(
        N_357), .Y(N_126));
    NOR2B DUMPTIME_1_sqmuxa (.A(top_code_0_pluseload), .B(
        top_code_0_pluse_lc), .Y(DUMPTIME_1_sqmuxa_net_1));
    MX2C \timecount_1_RNO_0[13]  (.A(\PLUSETIME[13]_net_1 ), .B(
        \DUMPTIME[13]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_100));
    AO1A off_test_RNO_0 (.A(\CS[5]_net_1 ), .B(plusestate_0_off_test), 
        .C(\CS[4]_net_1 ), .Y(N_145));
    MX2C \timecount_1_RNO_0[11]  (.A(\PLUSETIME[11]_net_1 ), .B(
        \DUMPTIME[11]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_98));
    DFN1 tetw_pluse (.D(N_61), .CLK(GLA), .Q(plusestate_0_tetw_pluse));
    AO1C \timecount_1_RNO[0]  (.A(N_153), .B(\PLUSETIME[0]_net_1 ), .C(
        \timecount_5_1_0[0] ), .Y(\timecount_5[0] ));
    OR2 \CS_RNIDRQ7[3]  (.A(\CS[4]_net_1 ), .B(\CS[3]_net_1 ), .Y(N_92)
        );
    MX2C \CS_RNO_0[9]  (.A(\CS[9]_net_1 ), .B(\CS[4]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_110));
    DFN1E1 \timecount_1[6]  (.D(N_15), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[6]));
    AO1C \timecount_1_RNO_1[7]  (.A(\DUMPTIME[7]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[7] ));
    NOR2 \timecount_1_RNO_2[3]  (.A(\PLUSETIME[3]_net_1 ), .B(N_153), 
        .Y(N_122));
    DFN1 \CS[7]  (.D(\CS_RNO[7]_net_1 ), .CLK(GLA), .Q(\CS[7]_net_1 ));
    NOR2 \timecount_1_RNO[15]  (.A(N_102), .B(N_71), .Y(N_33));
    DFN1 \CS[6]  (.D(\CS_RNO[6]_net_1 ), .CLK(GLA), .Q(\CS[6]_net_1 ));
    DFN1E1 \DUMPTIME[3]  (.D(plusedata[3]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[3]_net_1 ));
    DFN1 sw_acq1 (.D(N_151), .CLK(GLA), .Q(plusestate_0_sw_acq1));
    AO1B state_over_n_RNO (.A(plusestate_0_state_over_n), .B(N_354), 
        .C(top_code_0_pluse_rst), .Y(state_over_n_RNO_net_1));
    AOI1B \timecount_1_RNO_0[0]  (.A(\DUMPTIME[0]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_1_0[0] ));
    DFN1 dds_config (.D(N_57), .CLK(GLA), .Q(plusestate_0_dds_config));
    AO1C \timecount_1_RNO_1[3]  (.A(\DUMPTIME[3]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[3] ));
    OR2 \timecount_1_RNO_0[6]  (.A(\PLUSETIME[6]_net_1 ), .B(N_153), 
        .Y(N_135));
    NOR2A \CS_RNO[2]  (.A(top_code_0_pluse_rst_0), .B(N_104), .Y(
        \CS_RNO[2]_net_1 ));
    GND GND_i_0 (.Y(GND_0));
    DFN1 \CS[8]  (.D(\CS_RNO[8]_net_1 ), .CLK(GLA), .Q(\CS[8]_net_1 ));
    DFN1E1 \DUMPTIME[15]  (.D(plusedata[15]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[15]_net_1 ));
    MX2C \CS_RNO_0[8]  (.A(\CS[8]_net_1 ), .B(\CS[2]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_109));
    OR2 \timecount_1_RNO_0[8]  (.A(\PLUSETIME[8]_net_1 ), .B(N_153), 
        .Y(N_140));
    NOR3 \timecount_1_RNO[1]  (.A(N_116), .B(\timecount_5_i_0[1] ), .C(
        N_115), .Y(N_5));
    DFN1 pluse_acq (.D(N_63), .CLK(GLA), .Q(plusestate_0_pluse_acq));
    DFN1E1 \DUMPTIME[13]  (.D(plusedata[13]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[13]_net_1 ));
    NOR2 \CS_RNIJJR7[6]  (.A(\CS[7]_net_1 ), .B(\CS[6]_net_1 ), .Y(
        N_354));
    DFN1 \CS[2]  (.D(\CS_RNO[2]_net_1 ), .CLK(GLA), .Q(\CS[2]_net_1 ));
    OA1A \timecount_1_RNO_1[6]  (.A(\CS[5]_net_1 ), .B(
        \DUMPTIME[6]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[6] ));
    NOR2 \timecount_1_RNO_2[1]  (.A(\PLUSETIME[1]_net_1 ), .B(N_153), 
        .Y(N_115));
    OA1A tetw_pluse_RNO (.A(N_354), .B(plusestate_0_tetw_pluse), .C(
        top_code_0_pluse_rst_0), .Y(N_61));
    DFN1E1 \PLUSETIME[6]  (.D(plusedata[6]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[6]_net_1 ));
    DFN1E1 \PLUSETIME[13]  (.D(plusedata[13]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[13]_net_1 ));
    DFN1E1 \DUMPTIME[5]  (.D(plusedata[5]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[5]_net_1 ));
    NOR3A soft_d_RNO_1 (.A(N_354), .B(\CS[5]_net_1 ), .C(N_92), .Y(
        N_351));
    AO1C \timecount_1_RNO_1[1]  (.A(\DUMPTIME[1]_net_1 ), .B(
        \CS[5]_net_1 ), .C(top_code_0_pluse_rst_0), .Y(
        \timecount_5_i_0[1] ));
    NOR2 \timecount_1_RNO[13]  (.A(N_100), .B(N_71), .Y(N_29));
    NOR3A sw_acq1_RNO_1 (.A(N_354), .B(\CS[8]_net_1 ), .C(N_92), .Y(
        N_350));
    DFN1 off_test (.D(N_59), .CLK(GLA), .Q(plusestate_0_off_test));
    DFN1E1 \timecount_1[9]  (.D(N_21), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[9]));
    DFN1E1 \DUMPTIME[0]  (.D(plusedata[0]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[0]_net_1 ));
    NOR2B dds_config_RNO (.A(top_code_0_pluse_rst), .B(N_146), .Y(N_57)
        );
    DFN1E1 \PLUSETIME[0]  (.D(plusedata[0]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[0]_net_1 ));
    NOR2 \timecount_1_RNO[14]  (.A(N_101), .B(N_71), .Y(N_31));
    NOR2A \CS_RNO[8]  (.A(top_code_0_pluse_rst), .B(N_109), .Y(
        \CS_RNO[8]_net_1 ));
    DFN1 \CS[5]  (.D(\CS_RNO[5]_net_1 ), .CLK(GLA), .Q(\CS[5]_net_1 ));
    OA1B \timecount_1_RNO[2]  (.A(\CS[3]_net_1 ), .B(N_156), .C(
        \timecount_5_i_1[2] ), .Y(N_7));
    MX2C \CS_RNO_0[3]  (.A(\CS[3]_net_1 ), .B(\CS[8]_net_1 ), .S(
        timer_top_0_clk_en_pluse), .Y(N_105));
    DFN1E1 \PLUSETIME[2]  (.D(plusedata[2]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[2]_net_1 ));
    DFN1E1 \timecount_1[3]  (.D(N_9), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[3]));
    OR2 \CS_RNI9BQ7[1]  (.A(\CS[2]_net_1 ), .B(\CS[1]_net_1 ), .Y(N_91)
        );
    OR2 \CS_RNIKNR7_0[9]  (.A(\CS[9]_net_1 ), .B(\CS[5]_net_1 ), .Y(
        N_152));
    DFN1E1 \DUMPTIME[14]  (.D(plusedata[14]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[14]_net_1 ));
    DFN1E1 \DUMPTIME[11]  (.D(plusedata[11]), .CLK(GLA), .E(
        DUMPTIME_1_sqmuxa_net_1), .Q(\DUMPTIME[11]_net_1 ));
    NOR2 \timecount_1_RNO[9]  (.A(N_96), .B(N_71), .Y(N_21));
    DFN1E1 \PLUSETIME[7]  (.D(plusedata[7]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[7]_net_1 ));
    NOR2A \CS_RNO[6]  (.A(top_code_0_pluse_rst_0), .B(N_108), .Y(
        \CS_RNO[6]_net_1 ));
    OR2 \CS_RNIT2MF[1]  (.A(N_152), .B(N_91), .Y(N_156));
    NOR2 \timecount_1_RNO[11]  (.A(N_98), .B(N_71), .Y(N_25));
    OR2A \CS_RNI0G4E[6]  (.A(top_code_0_pluse_rst), .B(N_354), .Y(
        un1_sw_acq1_2_sqmuxa));
    AO1D \timecount_1_RNO_0[7]  (.A(\PLUSETIME[7]_net_1 ), .B(N_153), 
        .C(\timecount_5_i_0[7] ), .Y(\timecount_5_i_1[7] ));
    OR2 \CS_RNIFNPB[8]  (.A(N_152), .B(\CS[8]_net_1 ), .Y(N_155));
    NOR3C \timecount_1_RNO[8]  (.A(N_140), .B(\timecount_5_i_0[8] ), 
        .C(N_155), .Y(N_19));
    DFN1E1 \PLUSETIME[1]  (.D(plusedata[1]), .CLK(GLA), .E(
        DUMPTIME_0_sqmuxa_net_1), .Q(\PLUSETIME[1]_net_1 ));
    DFN1E1 \timecount_1[4]  (.D(N_11), .CLK(GLA), .E(
        un1_sw_acq1_2_sqmuxa), .Q(timecount_1_1[4]));
    MX2C \timecount_1_RNO_0[15]  (.A(\PLUSETIME[15]_net_1 ), .B(
        \DUMPTIME[15]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_102));
    MX2C \timecount_1_RNO_0[14]  (.A(\PLUSETIME[14]_net_1 ), .B(
        \DUMPTIME[14]_net_1 ), .S(\CS[5]_net_1 ), .Y(N_101));
    
endmodule


module bridge_div(
       scaleddsdiv,
       top_code_0_bridge_load,
       GLA,
       bri_dump_sw_0_reset_out,
       ddsclkout_c,
       clk_4f_en,
       pd_pulse_en_c
    );
input  [5:0] scaleddsdiv;
input  top_code_0_bridge_load;
input  GLA;
input  bri_dump_sw_0_reset_out;
input  ddsclkout_c;
output clk_4f_en;
input  pd_pulse_en_c;

    wire N_15, \count_RNITQSU3[1]_net_1 , \count_RNISQSU3[0]_net_1 , 
        N_7, \count_RNIVQSU3[3]_net_1 , \DWACT_FINC_E[0] , 
        \un1_count_NE_1[0] , \count[1]_net_1 , \dataall[1]_net_1 , 
        \un1_count_2_i[0] , \un1_count_NE_0[0] , \count[0]_net_1 , 
        \dataall[0]_net_1 , \un1_count_i_3[0] , \clear1_n17_NE_1[0] , 
        \datahalf[0]_net_1 , \clear1_n17_1_i[0] , \clear1_n17_NE_0[0] , 
        \count[3]_net_1 , \un1_count_i[0] , \un1_count_3_i[0] , 
        \clear1_n17_NE_i[0] , \clear1_n17_2_i[0] , clk_4f_1_sqmuxa, 
        \dataall_1[2] , CO1, \dataall_1[1] , CO0, \dataall_1[3] , 
        clk_4f_reg1_net_1, clk_4f_reg2_net_1, \dataall_1[0] , 
        clear1_n18, clk_4f_5, clk_4f_net_1, \count_RNIUQSU3[2]_net_1 , 
        \count[2]_net_1 , \count_RNI0RSU3[4]_net_1 , \count[4]_net_1 , 
        \count_RNI1RSU3[5]_net_1 , \count[5]_net_1 , 
        \datahalf[1]_net_1 , \datahalf[2]_net_1 , \dataall[2]_net_1 , 
        \dataall[3]_net_1 , \count_5[0] , \count_5[1] , \count_5[2] , 
        \count_5[3] , \count_5[4] , \count_5[5] , N_4, N_12, GND, VCC, 
        GND_0, VCC_0;
    
    DFN1C0 \count[5]  (.D(\count_5[5] ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(\count[5]_net_1 ));
    DFN1E0C0 clk_4f (.D(clk_4f_5), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .E(clk_4f_1_sqmuxa), .Q(clk_4f_net_1)
        );
    XOR2 count_5_I_24 (.A(N_4), .B(\count_RNI1RSU3[5]_net_1 ), .Y(
        \count_5[5] ));
    XNOR2 \datahalf_RNIOH29[1]  (.A(\datahalf[1]_net_1 ), .B(
        \count[1]_net_1 ), .Y(\clear1_n17_1_i[0] ));
    DFN1C0 \count[1]  (.D(\count_5[1] ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(\count[1]_net_1 ));
    DFN1E1 \datahalf[1]  (.D(scaleddsdiv[1]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\datahalf[1]_net_1 ));
    MAJ3 dataall_1_1_CO1 (.A(scaleddsdiv[4]), .B(CO0), .C(
        scaleddsdiv[1]), .Y(CO1));
    DFN1P0 \count[0]  (.D(\count_5[0] ), .CLK(ddsclkout_c), .PRE(
        bri_dump_sw_0_reset_out), .Q(\count[0]_net_1 ));
    AND3 count_5_I_23 (.A(\DWACT_FINC_E[0] ), .B(
        \count_RNIVQSU3[3]_net_1 ), .C(\count_RNI0RSU3[4]_net_1 ), .Y(
        N_4));
    NOR2A clk_4f_reg2_RNIV6JF (.A(clk_4f_reg1_net_1), .B(
        clk_4f_reg2_net_1), .Y(clk_4f_en));
    VCC VCC_i (.Y(VCC));
    NOR3C \count_RNISQSU3[0]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[0]_net_1 ), .Y(\count_RNISQSU3[0]_net_1 ));
    NOR2A \count_RNI14HK[3]  (.A(\un1_count_i_3[0] ), .B(
        \count[3]_net_1 ), .Y(\clear1_n17_NE_0[0] ));
    XNOR2 \dataall_RNISOPC[3]  (.A(\dataall[3]_net_1 ), .B(
        \count[3]_net_1 ), .Y(\un1_count_3_i[0] ));
    XA1A \dataall_RNIDRFQ[0]  (.A(\count[0]_net_1 ), .B(
        \dataall[0]_net_1 ), .C(\un1_count_i_3[0] ), .Y(
        \un1_count_NE_0[0] ));
    DFN1E1 \dataall[0]  (.D(\dataall_1[0] ), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\dataall[0]_net_1 ));
    DFN1C0 clk_4f_reg2 (.D(clk_4f_reg1_net_1), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(clk_4f_reg2_net_1));
    NOR2B dataall_1_1_ANB0 (.A(scaleddsdiv[3]), .B(scaleddsdiv[0]), .Y(
        CO0));
    DFN1E1 \dataall[2]  (.D(\dataall_1[2] ), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\dataall[2]_net_1 ));
    DFN1C0 clk_4f_reg1 (.D(clk_4f_net_1), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(clk_4f_reg1_net_1));
    DFN1C0 \count[2]  (.D(\count_5[2] ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(\count[2]_net_1 ));
    INV count_5_I_4 (.A(\count_RNISQSU3[0]_net_1 ), .Y(\count_5[0] ));
    NOR3C \datahalf_RNI9POF1[0]  (.A(\clear1_n17_NE_0[0] ), .B(
        \clear1_n17_2_i[0] ), .C(\clear1_n17_NE_1[0] ), .Y(
        \clear1_n17_NE_i[0] ));
    MAJ3 dataall_1_1_CO2 (.A(scaleddsdiv[5]), .B(CO1), .C(
        scaleddsdiv[2]), .Y(\dataall_1[3] ));
    OR2 \datahalf_RNI4VLG3[0]  (.A(\un1_count_i[0] ), .B(
        \clear1_n17_NE_i[0] ), .Y(clear1_n18));
    GND GND_i (.Y(GND));
    DFN1E1 \dataall[1]  (.D(\dataall_1[1] ), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\dataall[1]_net_1 ));
    XOR2 count_5_I_9 (.A(N_15), .B(\count_RNIUQSU3[2]_net_1 ), .Y(
        \count_5[2] ));
    NOR3C \count_RNIUQSU3[2]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[2]_net_1 ), .Y(\count_RNIUQSU3[2]_net_1 ));
    XNOR2 \dataall_RNIQOPC[2]  (.A(\dataall[2]_net_1 ), .B(
        \count[2]_net_1 ), .Y(\un1_count_2_i[0] ));
    DFN1E1 \datahalf[0]  (.D(scaleddsdiv[0]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\datahalf[0]_net_1 ));
    AND3 count_5_I_16 (.A(\count_RNISQSU3[0]_net_1 ), .B(
        \count_RNITQSU3[1]_net_1 ), .C(\count_RNIUQSU3[2]_net_1 ), .Y(
        \DWACT_FINC_E[0] ));
    OR3C \dataall_RNIR5T02[0]  (.A(\un1_count_NE_0[0] ), .B(
        \un1_count_3_i[0] ), .C(\un1_count_NE_1[0] ), .Y(
        \un1_count_i[0] ));
    NOR2 \count_RNIN2MD[4]  (.A(\count[5]_net_1 ), .B(\count[4]_net_1 )
        , .Y(\un1_count_i_3[0] ));
    NOR2B count_5_I_8 (.A(\count_RNITQSU3[1]_net_1 ), .B(
        \count_RNISQSU3[0]_net_1 ), .Y(N_15));
    XOR2 count_5_I_5 (.A(\count_RNISQSU3[0]_net_1 ), .B(
        \count_RNITQSU3[1]_net_1 ), .Y(\count_5[1] ));
    XA1A \datahalf_RNIEV4I[0]  (.A(\count[0]_net_1 ), .B(
        \datahalf[0]_net_1 ), .C(\clear1_n17_1_i[0] ), .Y(
        \clear1_n17_NE_1[0] ));
    XOR3 dataall_1_1_SUM2_0 (.A(scaleddsdiv[2]), .B(scaleddsdiv[5]), 
        .C(CO1), .Y(\dataall_1[2] ));
    NOR3C \count_RNITQSU3[1]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[1]_net_1 ), .Y(\count_RNITQSU3[1]_net_1 ));
    NOR3C \count_RNIVQSU3[3]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[3]_net_1 ), .Y(\count_RNIVQSU3[3]_net_1 ));
    DFN1C0 \count[3]  (.D(\count_5[3] ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(\count[3]_net_1 ));
    NOR3C \count_RNI1RSU3[5]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[5]_net_1 ), .Y(\count_RNI1RSU3[5]_net_1 ));
    NOR2A clk_4f_RNO (.A(pd_pulse_en_c), .B(clk_4f_net_1), .Y(clk_4f_5)
        );
    XOR2 dataall_1_1_SUM0_0 (.A(scaleddsdiv[3]), .B(scaleddsdiv[0]), 
        .Y(\dataall_1[0] ));
    NOR2B count_5_I_19 (.A(\count_RNIVQSU3[3]_net_1 ), .B(
        \DWACT_FINC_E[0] ), .Y(N_7));
    XNOR2 \datahalf_RNIQL29[2]  (.A(\datahalf[2]_net_1 ), .B(
        \count[2]_net_1 ), .Y(\clear1_n17_2_i[0] ));
    DFN1E1 \datahalf[2]  (.D(scaleddsdiv[2]), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\datahalf[2]_net_1 ));
    NOR3B clk_4f_RNO_0 (.A(pd_pulse_en_c), .B(\un1_count_i[0] ), .C(
        \clear1_n17_NE_i[0] ), .Y(clk_4f_1_sqmuxa));
    DFN1E1 \dataall[3]  (.D(\dataall_1[3] ), .CLK(GLA), .E(
        top_code_0_bridge_load), .Q(\dataall[3]_net_1 ));
    XOR2 count_5_I_20 (.A(N_7), .B(\count_RNI0RSU3[4]_net_1 ), .Y(
        \count_5[4] ));
    XOR2 count_5_I_13 (.A(N_12), .B(\count_RNIVQSU3[3]_net_1 ), .Y(
        \count_5[3] ));
    DFN1C0 \count[4]  (.D(\count_5[4] ), .CLK(ddsclkout_c), .CLR(
        bri_dump_sw_0_reset_out), .Q(\count[4]_net_1 ));
    AND3 count_5_I_12 (.A(\count_RNISQSU3[0]_net_1 ), .B(
        \count_RNITQSU3[1]_net_1 ), .C(\count_RNIUQSU3[2]_net_1 ), .Y(
        N_12));
    XA1A \dataall_RNIIHJP[1]  (.A(\count[1]_net_1 ), .B(
        \dataall[1]_net_1 ), .C(\un1_count_2_i[0] ), .Y(
        \un1_count_NE_1[0] ));
    XOR3 dataall_1_1_SUM1_0 (.A(scaleddsdiv[1]), .B(scaleddsdiv[4]), 
        .C(CO0), .Y(\dataall_1[1] ));
    NOR3C \count_RNI0RSU3[4]  (.A(clear1_n18), .B(pd_pulse_en_c), .C(
        \count[4]_net_1 ), .Y(\count_RNI0RSU3[4]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module s_acq_change(
       s_acqnum_1,
       s_acqnum_0,
       strippluse,
       change,
       s_acqnum,
       s_stripnum,
       un1_top_code_0_3_0,
       s_acq_change_0_s_load,
       scalestate_0_load_out,
       top_code_0_s_load,
       net_45,
       net_33_0,
       net_27,
       s_acq_change_0_s_rst,
       GLA,
       s_acq_change_0_s_load_0
    );
input  [11:0] s_acqnum_1;
input  [15:0] s_acqnum_0;
input  [11:0] strippluse;
input  [1:0] change;
output [15:0] s_acqnum;
output [11:0] s_stripnum;
input  [1:0] un1_top_code_0_3_0;
output s_acq_change_0_s_load;
input  scalestate_0_load_out;
input  top_code_0_s_load;
input  net_45;
input  net_33_0;
input  net_27;
output s_acq_change_0_s_rst;
input  GLA;
output s_acq_change_0_s_load_0;

    wire s_load_0_0_RNIMC0R_net_1, s_rst_net_1, N_65, s_rst_5, N_66, 
        s_load_5_net_1, N_53, \s_stripnum_5[0] , N_54, 
        \s_stripnum_5[1] , N_55, \s_stripnum_5[2] , N_57, 
        \s_stripnum_5[4] , N_58, \s_stripnum_5[5] , N_59, 
        \s_stripnum_5[6] , N_60, \s_stripnum_5[7] , N_61, 
        \s_stripnum_5[8] , N_62, \s_stripnum_5[9] , N_63, 
        \s_stripnum_5[10] , N_64, \s_stripnum_5[11] , N_67, 
        \s_acqnum_5[0] , N_68, \s_acqnum_5[1] , N_69, \s_acqnum_5[2] , 
        N_70, \s_acqnum_5[3] , N_71, \s_acqnum_5[4] , N_72, 
        \s_acqnum_5[5] , N_73, \s_acqnum_5[6] , N_74, \s_acqnum_5[7] , 
        N_75, \s_acqnum_5[8] , N_77, \s_acqnum_5[10] , N_78, 
        \s_acqnum_5[11] , N_79, \s_acqnum_5[12] , N_80, 
        \s_acqnum_5[13] , N_81, \s_acqnum_5[14] , N_82, 
        \s_acqnum_5[15] , s_rst_RNO_net_1, \s_stripnum_RNO[0]_net_1 , 
        \s_stripnum_RNO[1]_net_1 , \s_acqnum_RNO[3]_net_1 , 
        \s_acqnum_RNO[4]_net_1 , \s_acqnum_RNO[5]_net_1 , 
        \s_acqnum_RNO[6]_net_1 , \s_acqnum_RNO[7]_net_1 , 
        \s_acqnum_RNO[8]_net_1 , \s_acqnum_RNO[10]_net_1 , 
        \s_acqnum_RNO[11]_net_1 , \s_acqnum_RNO[12]_net_1 , 
        \s_acqnum_RNO[13]_net_1 , \s_acqnum_RNO[14]_net_1 , 
        \s_acqnum_RNO[15]_net_1 , \s_stripnum_RNO[2]_net_1 , 
        \s_stripnum_RNO[4]_net_1 , \s_stripnum_RNO[5]_net_1 , 
        \s_stripnum_RNO[6]_net_1 , \s_stripnum_RNO[7]_net_1 , 
        \s_stripnum_RNO[8]_net_1 , \s_stripnum_RNO[9]_net_1 , 
        \s_stripnum_RNO[10]_net_1 , \s_stripnum_RNO[11]_net_1 , 
        \s_acqnum_RNO[0]_net_1 , \s_acqnum_RNO[1]_net_1 , 
        \s_acqnum_RNO[2]_net_1 , \s_stripnum_5[3] , \s_acqnum_5[9] , 
        \s_stripnum_RNO[3]_net_1 , N_56, \s_acqnum_RNO[9]_net_1 , N_76, 
        GND, VCC, GND_0, VCC_0;
    
    DFN1 \s_stripnum[4]  (.D(\s_stripnum_RNO[4]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[4]));
    DFN1 s_load (.D(s_load_0_0_RNIMC0R_net_1), .CLK(GLA), .Q(
        s_acq_change_0_s_load));
    MX2 \s_acqnum_RNO_0[13]  (.A(\s_acqnum_5[13] ), .B(s_acqnum[13]), 
        .S(change[1]), .Y(N_80));
    NOR2B \s_stripnum_RNO_1[2]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[2]), .Y(\s_stripnum_5[2] ));
    NOR2B \s_stripnum_RNO[7]  (.A(N_60), .B(net_27), .Y(
        \s_stripnum_RNO[7]_net_1 ));
    NOR2A \s_acqnum_RNO_1[13]  (.A(s_acqnum_0[13]), .B(change[0]), .Y(
        \s_acqnum_5[13] ));
    NOR2B \s_acqnum_RNO[14]  (.A(N_81), .B(net_27), .Y(
        \s_acqnum_RNO[14]_net_1 ));
    NOR2B s_rst_RNO (.A(N_65), .B(net_27), .Y(s_rst_RNO_net_1));
    NOR2B \s_stripnum_RNO_1[8]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[8]), .Y(\s_stripnum_5[8] ));
    DFN1 \s_acqnum[9]  (.D(\s_acqnum_RNO[9]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[9]));
    NOR2B \s_stripnum_RNO_1[1]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[1]), .Y(\s_stripnum_5[1] ));
    NOR2B \s_stripnum_RNO_1[9]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[9]), .Y(\s_stripnum_5[9] ));
    DFN1 \s_stripnum[1]  (.D(\s_stripnum_RNO[1]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[1]));
    MX2 \s_acqnum_RNO_0[7]  (.A(\s_acqnum_5[7] ), .B(s_acqnum[7]), .S(
        change[1]), .Y(N_74));
    MX2 \s_acqnum_RNO_0[14]  (.A(\s_acqnum_5[14] ), .B(s_acqnum[14]), 
        .S(change[1]), .Y(N_81));
    NOR2A \s_acqnum_RNO_1[14]  (.A(s_acqnum_0[14]), .B(change[0]), .Y(
        \s_acqnum_5[14] ));
    MX2 \s_stripnum_RNO_0[2]  (.A(\s_stripnum_5[2] ), .B(s_stripnum[2])
        , .S(un1_top_code_0_3_0[1]), .Y(N_55));
    NOR2B \s_stripnum_RNO_1[10]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[10]), .Y(\s_stripnum_5[10] ));
    MX2 s_load_0_0_RNIUU5P (.A(s_load_5_net_1), .B(
        s_acq_change_0_s_load_0), .S(un1_top_code_0_3_0[1]), .Y(N_66));
    DFN1 \s_acqnum[2]  (.D(\s_acqnum_RNO[2]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[2]));
    VCC VCC_i (.Y(VCC));
    NOR2B \s_stripnum_RNO_1[11]  (.A(change[0]), .B(strippluse[11]), 
        .Y(\s_stripnum_5[11] ));
    NOR2B \s_stripnum_RNO[11]  (.A(N_64), .B(net_27), .Y(
        \s_stripnum_RNO[11]_net_1 ));
    NOR2B \s_stripnum_RNO_1[5]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[5]), .Y(\s_stripnum_5[5] ));
    NOR2B \s_stripnum_RNO[2]  (.A(N_55), .B(net_27), .Y(
        \s_stripnum_RNO[2]_net_1 ));
    MX2 s_load_5 (.A(top_code_0_s_load), .B(scalestate_0_load_out), .S(
        change[0]), .Y(s_load_5_net_1));
    MX2 \s_stripnum_RNO_0[5]  (.A(\s_stripnum_5[5] ), .B(s_stripnum[5])
        , .S(un1_top_code_0_3_0[1]), .Y(N_58));
    CLKINT s_rst_RNI2O37 (.A(s_rst_net_1), .Y(s_acq_change_0_s_rst));
    NOR2B \s_acqnum_RNO[15]  (.A(N_82), .B(net_27), .Y(
        \s_acqnum_RNO[15]_net_1 ));
    NOR2B \s_stripnum_RNO_1[3]  (.A(change[0]), .B(strippluse[3]), .Y(
        \s_stripnum_5[3] ));
    NOR2B \s_acqnum_RNO[3]  (.A(N_70), .B(net_27), .Y(
        \s_acqnum_RNO[3]_net_1 ));
    MX2 \s_acqnum_RNO_1[3]  (.A(s_acqnum_0[3]), .B(s_acqnum_1[3]), .S(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[3] ));
    NOR2B \s_acqnum_RNO[0]  (.A(N_67), .B(net_27), .Y(
        \s_acqnum_RNO[0]_net_1 ));
    MX2 \s_acqnum_RNO_1[5]  (.A(s_acqnum_0[5]), .B(s_acqnum_1[5]), .S(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[5] ));
    MX2 \s_acqnum_RNO_0[1]  (.A(\s_acqnum_5[1] ), .B(s_acqnum[1]), .S(
        un1_top_code_0_3_0[1]), .Y(N_68));
    DFN1 \s_stripnum[9]  (.D(\s_stripnum_RNO[9]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[9]));
    DFN1 \s_stripnum[6]  (.D(\s_stripnum_RNO[6]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[6]));
    NOR2B \s_stripnum_RNO[5]  (.A(N_58), .B(net_27), .Y(
        \s_stripnum_RNO[5]_net_1 ));
    DFN1 s_rst (.D(s_rst_RNO_net_1), .CLK(GLA), .Q(s_rst_net_1));
    MX2 \s_acqnum_RNO_1[7]  (.A(s_acqnum_0[7]), .B(s_acqnum_1[7]), .S(
        change[0]), .Y(\s_acqnum_5[7] ));
    NOR2B \s_stripnum_RNO[4]  (.A(N_57), .B(net_27), .Y(
        \s_stripnum_RNO[4]_net_1 ));
    DFN1 \s_acqnum[4]  (.D(\s_acqnum_RNO[4]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[4]));
    DFN1 \s_acqnum[8]  (.D(\s_acqnum_RNO[8]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[8]));
    MX2 \s_stripnum_RNO_0[7]  (.A(\s_stripnum_5[7] ), .B(s_stripnum[7])
        , .S(un1_top_code_0_3_0[1]), .Y(N_60));
    MX2 \s_acqnum_RNO_0[5]  (.A(\s_acqnum_5[5] ), .B(s_acqnum[5]), .S(
        change[1]), .Y(N_72));
    DFN1 \s_stripnum[3]  (.D(\s_stripnum_RNO[3]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[3]));
    MX2 \s_acqnum_RNO_1[0]  (.A(s_acqnum_0[0]), .B(s_acqnum_1[0]), .S(
        change[0]), .Y(\s_acqnum_5[0] ));
    NOR2B \s_acqnum_RNO[5]  (.A(N_72), .B(net_27), .Y(
        \s_acqnum_RNO[5]_net_1 ));
    NOR2B \s_acqnum_RNO[2]  (.A(N_69), .B(net_27), .Y(
        \s_acqnum_RNO[2]_net_1 ));
    MX2 \s_acqnum_RNO_0[10]  (.A(\s_acqnum_5[10] ), .B(s_acqnum[10]), 
        .S(change[1]), .Y(N_77));
    MX2 \s_stripnum_RNO_0[6]  (.A(\s_stripnum_5[6] ), .B(s_stripnum[6])
        , .S(un1_top_code_0_3_0[1]), .Y(N_59));
    MX2 \s_acqnum_RNO_1[10]  (.A(s_acqnum_0[10]), .B(s_acqnum_1[10]), 
        .S(un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[10] ));
    MX2 \s_stripnum_RNO_0[1]  (.A(\s_stripnum_5[1] ), .B(s_stripnum[1])
        , .S(un1_top_code_0_3_0[1]), .Y(N_54));
    MX2 \s_acqnum_RNO_0[8]  (.A(\s_acqnum_5[8] ), .B(s_acqnum[8]), .S(
        change[1]), .Y(N_75));
    DFN1 \s_acqnum[12]  (.D(\s_acqnum_RNO[12]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[12]));
    NOR2B \s_stripnum_RNO[8]  (.A(N_61), .B(net_27), .Y(
        \s_stripnum_RNO[8]_net_1 ));
    DFN1 \s_acqnum[1]  (.D(\s_acqnum_RNO[1]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[1]));
    DFN1 \s_acqnum[15]  (.D(\s_acqnum_RNO[15]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[15]));
    NOR2B \s_acqnum_RNO[11]  (.A(N_78), .B(net_27), .Y(
        \s_acqnum_RNO[11]_net_1 ));
    DFN1 \s_acqnum[11]  (.D(\s_acqnum_RNO[11]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[11]));
    NOR2B \s_acqnum_RNO[12]  (.A(N_79), .B(net_27), .Y(
        \s_acqnum_RNO[12]_net_1 ));
    DFN1 \s_acqnum[7]  (.D(\s_acqnum_RNO[7]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[7]));
    DFN1 \s_acqnum[0]  (.D(\s_acqnum_RNO[0]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[0]));
    GND GND_i (.Y(GND));
    MX2 \s_stripnum_RNO_0[10]  (.A(\s_stripnum_5[10] ), .B(
        s_stripnum[10]), .S(un1_top_code_0_3_0[1]), .Y(N_63));
    NOR2B \s_stripnum_RNO[0]  (.A(N_53), .B(net_27), .Y(
        \s_stripnum_RNO[0]_net_1 ));
    MX2 \s_acqnum_RNO_1[6]  (.A(s_acqnum_0[6]), .B(s_acqnum_1[6]), .S(
        change[0]), .Y(\s_acqnum_5[6] ));
    MX2 \s_acqnum_RNO_0[3]  (.A(\s_acqnum_5[3] ), .B(s_acqnum[3]), .S(
        un1_top_code_0_3_0[1]), .Y(N_70));
    DFN1 \s_stripnum[5]  (.D(\s_stripnum_RNO[5]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[5]));
    MX2 \s_stripnum_RNO_0[11]  (.A(\s_stripnum_5[11] ), .B(
        s_stripnum[11]), .S(un1_top_code_0_3_0[1]), .Y(N_64));
    NOR2B \s_acqnum_RNO[4]  (.A(N_71), .B(net_27), .Y(
        \s_acqnum_RNO[4]_net_1 ));
    NOR2B \s_stripnum_RNO[3]  (.A(N_56), .B(net_27), .Y(
        \s_stripnum_RNO[3]_net_1 ));
    NOR2B s_load_0_0_RNIMC0R (.A(N_66), .B(net_27), .Y(
        s_load_0_0_RNIMC0R_net_1));
    NOR2B \s_acqnum_RNO[13]  (.A(N_80), .B(net_27), .Y(
        \s_acqnum_RNO[13]_net_1 ));
    NOR2B \s_stripnum_RNO_1[6]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[6]), .Y(\s_stripnum_5[6] ));
    MX2 \s_acqnum_RNO_0[9]  (.A(\s_acqnum_5[9] ), .B(s_acqnum[9]), .S(
        change[1]), .Y(N_76));
    NOR2B \s_acqnum_RNO[8]  (.A(N_75), .B(net_27), .Y(
        \s_acqnum_RNO[8]_net_1 ));
    NOR2B \s_stripnum_RNO[9]  (.A(N_62), .B(net_27), .Y(
        \s_stripnum_RNO[9]_net_1 ));
    DFN1 \s_stripnum[11]  (.D(\s_stripnum_RNO[11]_net_1 ), .CLK(GLA), 
        .Q(s_stripnum[11]));
    DFN1 \s_acqnum[14]  (.D(\s_acqnum_RNO[14]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[14]));
    NOR2B \s_stripnum_RNO[6]  (.A(N_59), .B(net_27), .Y(
        \s_stripnum_RNO[6]_net_1 ));
    MX2 \s_acqnum_RNO_1[4]  (.A(s_acqnum_0[4]), .B(s_acqnum_1[4]), .S(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[4] ));
    DFN1 \s_stripnum[10]  (.D(\s_stripnum_RNO[10]_net_1 ), .CLK(GLA), 
        .Q(s_stripnum[10]));
    MX2 \s_acqnum_RNO_1[9]  (.A(s_acqnum_0[9]), .B(s_acqnum_1[9]), .S(
        change[0]), .Y(\s_acqnum_5[9] ));
    DFN1 \s_stripnum[7]  (.D(\s_stripnum_RNO[7]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[7]));
    MX2 \s_acqnum_RNO_1[8]  (.A(s_acqnum_0[8]), .B(s_acqnum_1[8]), .S(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[8] ));
    DFN1 \s_acqnum[6]  (.D(\s_acqnum_RNO[6]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[6]));
    NOR2B \s_acqnum_RNO[1]  (.A(N_68), .B(net_27), .Y(
        \s_acqnum_RNO[1]_net_1 ));
    MX2 \s_stripnum_RNO_0[4]  (.A(\s_stripnum_5[4] ), .B(s_stripnum[4])
        , .S(un1_top_code_0_3_0[1]), .Y(N_57));
    NOR2B \s_stripnum_RNO[10]  (.A(N_63), .B(net_27), .Y(
        \s_stripnum_RNO[10]_net_1 ));
    NOR2B \s_stripnum_RNO_1[7]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[7]), .Y(\s_stripnum_5[7] ));
    DFN1 \s_acqnum[10]  (.D(\s_acqnum_RNO[10]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[10]));
    NOR2B \s_stripnum_RNO_1[4]  (.A(un1_top_code_0_3_0[0]), .B(
        strippluse[4]), .Y(\s_stripnum_5[4] ));
    NOR2B \s_stripnum_RNO_1[0]  (.A(change[0]), .B(strippluse[0]), .Y(
        \s_stripnum_5[0] ));
    DFN1 \s_stripnum[8]  (.D(\s_stripnum_RNO[8]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[8]));
    DFN1 \s_stripnum[2]  (.D(\s_stripnum_RNO[2]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[2]));
    MX2 \s_acqnum_RNO_1[2]  (.A(s_acqnum_0[2]), .B(s_acqnum_1[2]), .S(
        change[0]), .Y(\s_acqnum_5[2] ));
    NOR2B \s_acqnum_RNO[10]  (.A(N_77), .B(net_27), .Y(
        \s_acqnum_RNO[10]_net_1 ));
    DFN1 \s_acqnum[5]  (.D(\s_acqnum_RNO[5]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[5]));
    DFN1 \s_acqnum[13]  (.D(\s_acqnum_RNO[13]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[13]));
    MX2 \s_stripnum_RNO_0[3]  (.A(\s_stripnum_5[3] ), .B(s_stripnum[3])
        , .S(change[1]), .Y(N_56));
    MX2 \s_stripnum_RNO_0[0]  (.A(\s_stripnum_5[0] ), .B(s_stripnum[0])
        , .S(un1_top_code_0_3_0[1]), .Y(N_53));
    MX2 \s_acqnum_RNO_1[1]  (.A(s_acqnum_0[1]), .B(s_acqnum_1[1]), .S(
        change[0]), .Y(\s_acqnum_5[1] ));
    MX2 \s_acqnum_RNO_0[0]  (.A(\s_acqnum_5[0] ), .B(s_acqnum[0]), .S(
        un1_top_code_0_3_0[1]), .Y(N_67));
    NOR2B \s_acqnum_RNO[6]  (.A(N_73), .B(net_27), .Y(
        \s_acqnum_RNO[6]_net_1 ));
    MX2 \s_acqnum_RNO_0[4]  (.A(\s_acqnum_5[4] ), .B(s_acqnum[4]), .S(
        change[1]), .Y(N_71));
    MX2 \s_acqnum_RNO_0[6]  (.A(\s_acqnum_5[6] ), .B(s_acqnum[6]), .S(
        change[1]), .Y(N_73));
    DFN1 \s_acqnum[3]  (.D(\s_acqnum_RNO[3]_net_1 ), .CLK(GLA), .Q(
        s_acqnum[3]));
    NOR2B \s_stripnum_RNO[1]  (.A(N_54), .B(net_27), .Y(
        \s_stripnum_RNO[1]_net_1 ));
    MX2 \s_acqnum_RNO_0[15]  (.A(\s_acqnum_5[15] ), .B(s_acqnum[15]), 
        .S(change[1]), .Y(N_82));
    NOR2A \s_acqnum_RNO_1[15]  (.A(s_acqnum_0[15]), .B(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[15] ));
    MX2 \s_acqnum_RNO_0[11]  (.A(\s_acqnum_5[11] ), .B(s_acqnum[11]), 
        .S(change[1]), .Y(N_78));
    NOR2B \s_acqnum_RNO[9]  (.A(N_76), .B(net_27), .Y(
        \s_acqnum_RNO[9]_net_1 ));
    MX2 s_rst_RNO_0 (.A(s_rst_5), .B(s_acq_change_0_s_rst), .S(
        un1_top_code_0_3_0[1]), .Y(N_65));
    MX2 \s_acqnum_RNO_1[11]  (.A(s_acqnum_0[11]), .B(s_acqnum_1[11]), 
        .S(un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[11] ));
    DFN1 s_load_0_0 (.D(s_load_0_0_RNIMC0R_net_1), .CLK(GLA), .Q(
        s_acq_change_0_s_load_0));
    NOR2B \s_acqnum_RNO[7]  (.A(N_74), .B(net_27), .Y(
        \s_acqnum_RNO[7]_net_1 ));
    DFN1 \s_stripnum[0]  (.D(\s_stripnum_RNO[0]_net_1 ), .CLK(GLA), .Q(
        s_stripnum[0]));
    MX2 \s_stripnum_RNO_0[8]  (.A(\s_stripnum_5[8] ), .B(s_stripnum[8])
        , .S(un1_top_code_0_3_0[1]), .Y(N_61));
    MX2 \s_acqnum_RNO_0[2]  (.A(\s_acqnum_5[2] ), .B(s_acqnum[2]), .S(
        un1_top_code_0_3_0[1]), .Y(N_69));
    MX2 \s_acqnum_RNO_0[12]  (.A(\s_acqnum_5[12] ), .B(s_acqnum[12]), 
        .S(change[1]), .Y(N_79));
    MX2 \s_stripnum_RNO_0[9]  (.A(\s_stripnum_5[9] ), .B(s_stripnum[9])
        , .S(un1_top_code_0_3_0[1]), .Y(N_62));
    NOR2A \s_acqnum_RNO_1[12]  (.A(s_acqnum_0[12]), .B(
        un1_top_code_0_3_0[0]), .Y(\s_acqnum_5[12] ));
    VCC VCC_i_0 (.Y(VCC_0));
    MX2 s_rst_RNO_1 (.A(net_33_0), .B(net_45), .S(change[0]), .Y(
        s_rst_5));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_3(
       count_9,
       GLA,
       state1ms_choice_0_reset_out,
       dump_state_0_off_start,
       off_on_state_0_state_over
    );
output [4:0] count_9;
input  GLA;
input  state1ms_choice_0_reset_out;
input  dump_state_0_off_start;
input  off_on_state_0_state_over;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_14, GND, VCC, GND_0, VCC_0;
    
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_9[0]), .B(count_9[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_9[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_9[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count_9[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    NOR2B \count_RNO_0[4]  (.A(count_9[3]), .B(N_13), .Y(N_14));
    NOR2B \count_RNIDKTJ[2]  (.A(count_9[2]), .B(N_12), .Y(N_13));
    XA1B \count_RNO[2]  (.A(N_12), .B(count_9[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(off_on_state_0_state_over), .B(
        dump_state_0_off_start), .C(state1ms_choice_0_reset_out), .Y(
        count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2B \count_RNITU8D[1]  (.A(count_9[1]), .B(count_9[0]), .Y(N_12));
    XA1B \count_RNO[4]  (.A(N_14), .B(count_9[4]), .C(
        count_0_sqmuxa_net_1), .Y(N_11));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_9[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_9[4]));
    NOR2 \count_RNO[0]  (.A(count_9[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_9[2]));
    
endmodule


module dump_state(
       i_9,
       i_8,
       i_5,
       i_1,
       i_0,
       dump_state_0_off_start,
       GLA,
       state1ms_choice_0_reset_out,
       dump_state_0_timer_start,
       dump_state_0_on_start
    );
input  [0:0] i_9;
input  [1:1] i_8;
input  [3:2] i_5;
input  [5:4] i_1;
input  [8:6] i_0;
output dump_state_0_off_start;
input  GLA;
input  state1ms_choice_0_reset_out;
output dump_state_0_timer_start;
output dump_state_0_on_start;

    wire un1_ns_0_a3_0, N_206_i, N_201, \cs_RNO_4[5] , cs4, N_193, 
        \cs_RNO_1[5]_net_1 , N_167, \cs[6]_net_1 , N_203, 
        \cs_RNO_3[4] , N_185, N_186, \cs_RNO_2[2] , N_182, N_183, 
        \cs[4]_net_1 , \cs_nsss[6] , N_166, N_2026_tz_tz, N_88, N_168, 
        \ns[3] , \cs_nsss_i[1] , N_171, \cs[1]_net_1 , \cs[2]_net_1 , 
        \cs_nsss[3] , N_195, N_196, \cs[3]_net_1 , N_173, \cs_nsss[7] , 
        off_start_RNO_net_1, N_176, \cs[7]_net_1 , \cs_i_0[0]_net_1 , 
        timer_start_RNO_net_1, GND, VCC, GND_0, VCC_0;
    
    DFN1 off_start (.D(off_start_RNO_net_1), .CLK(GLA), .Q(
        dump_state_0_off_start));
    NOR2B \cs_RNO_3[5]  (.A(i_5[3]), .B(\cs[4]_net_1 ), .Y(
        N_2026_tz_tz));
    DFN1 timer_start (.D(timer_start_RNO_net_1), .CLK(GLA), .Q(
        dump_state_0_timer_start));
    AO1B timer_start_RNO_0 (.A(dump_state_0_timer_start), .B(N_168), 
        .C(\ns[3] ), .Y(N_88));
    DFN1 \cs[6]  (.D(\cs_nsss[6] ), .CLK(GLA), .Q(\cs[6]_net_1 ));
    OR2A \cs_RNIHCFG[5]  (.A(dump_state_0_on_start), .B(N_206_i), .Y(
        un1_ns_0_a3_0));
    AO1C \cs_i_0_RNIIHUB[0]  (.A(i_8[1]), .B(\cs[1]_net_1 ), .C(
        \cs_i_0[0]_net_1 ), .Y(N_171));
    NOR2B timer_start_RNO (.A(cs4), .B(N_88), .Y(timer_start_RNO_net_1)
        );
    VCC VCC_i (.Y(VCC));
    DFN1 \cs[3]  (.D(\cs_nsss[3] ), .CLK(GLA), .Q(\cs[3]_net_1 ));
    NOR2A \cs_RNO[7]  (.A(cs4), .B(N_168), .Y(\cs_nsss[7] ));
    NOR2B \cs_RNO[1]  (.A(cs4), .B(N_171), .Y(\cs_nsss_i[1] ));
    DFN1 \cs[5]  (.D(\cs_RNO_4[5] ), .CLK(GLA), .Q(
        dump_state_0_on_start));
    DFN1 \cs_i_0[0]  (.D(cs4), .CLK(GLA), .Q(\cs_i_0[0]_net_1 ));
    NOR2B \cs_RNI5KH9[3]  (.A(i_8[1]), .B(\cs[3]_net_1 ), .Y(N_195));
    OA1C timer_start_RNO_1 (.A(\cs[3]_net_1 ), .B(i_8[1]), .C(N_173), 
        .Y(\ns[3] ));
    OR3A un1_ns_0_a2 (.A(i_0[8]), .B(i_1[4]), .C(i_0[6]), .Y(N_201));
    AO1A off_start_RNO (.A(N_176), .B(cs4), .C(\cs_nsss[6] ), .Y(
        off_start_RNO_net_1));
    DFN1 \cs[2]  (.D(\cs_RNO_2[2] ), .CLK(GLA), .Q(\cs[2]_net_1 ));
    NOR2B \cs_RNI5OH9[2]  (.A(i_5[2]), .B(\cs[2]_net_1 ), .Y(N_196));
    GND GND_i (.Y(GND));
    NOR3 off_start_RNO_0 (.A(N_195), .B(N_196), .C(N_171), .Y(N_176));
    AOI1 \cs_RNIUK1Q[6]  (.A(dump_state_0_on_start), .B(N_203), .C(
        \cs[6]_net_1 ), .Y(N_166));
    NOR3A \cs_RNO[2]  (.A(cs4), .B(N_182), .C(N_183), .Y(\cs_RNO_2[2] )
        );
    OA1B \cs_RNI9TR71[7]  (.A(N_201), .B(un1_ns_0_a3_0), .C(
        \cs[7]_net_1 ), .Y(N_168));
    NOR2A \cs_RNO_1[4]  (.A(i_8[1]), .B(\cs[4]_net_1 ), .Y(N_186));
    AOI1 \cs_RNO_0[2]  (.A(i_8[1]), .B(\cs[1]_net_1 ), .C(
        \cs[2]_net_1 ), .Y(N_182));
    NOR3 \cs_RNO_1[5]  (.A(dump_state_0_on_start), .B(\cs[6]_net_1 ), 
        .C(N_2026_tz_tz), .Y(\cs_RNO_1[5]_net_1 ));
    NOR2A \cs_RNI8SH9[4]  (.A(\cs[4]_net_1 ), .B(i_5[3]), .Y(N_173));
    NOR2B cs4_0_o3 (.A(state1ms_choice_0_reset_out), .B(i_9[0]), .Y(
        cs4));
    NOR3A \cs_RNO[4]  (.A(cs4), .B(N_185), .C(N_186), .Y(\cs_RNO_3[4] )
        );
    OR2 \cs_srsts_0_0_a2_0[6]  (.A(i_0[7]), .B(i_1[5]), .Y(N_206_i));
    NOR3 \cs_RNO_0[5]  (.A(N_206_i), .B(\cs[4]_net_1 ), .C(N_167), .Y(
        N_193));
    NOR3A \cs_RNI68PG1[6]  (.A(cs4), .B(N_166), .C(N_206_i), .Y(
        \cs_nsss[6] ));
    NOR2A \cs_RNO_1[2]  (.A(i_5[2]), .B(\cs[1]_net_1 ), .Y(N_183));
    NOR3A \cs_RNO_2[5]  (.A(N_201), .B(\cs[6]_net_1 ), .C(N_203), .Y(
        N_167));
    XA1B \cs_srsts_0_0_a2_1[6]  (.A(i_1[4]), .B(i_0[6]), .C(i_0[8]), 
        .Y(N_203));
    OA1 \cs_RNO[3]  (.A(N_195), .B(N_196), .C(cs4), .Y(\cs_nsss[3] ));
    DFN1 \cs[1]  (.D(\cs_nsss_i[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    NOR3A \cs_RNO[5]  (.A(cs4), .B(N_193), .C(\cs_RNO_1[5]_net_1 ), .Y(
        \cs_RNO_4[5] ));
    DFN1 \cs[4]  (.D(\cs_RNO_3[4] ), .CLK(GLA), .Q(\cs[4]_net_1 ));
    DFN1 \cs[7]  (.D(\cs_nsss[7] ), .CLK(GLA), .Q(\cs[7]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR2 \cs_RNO_0[4]  (.A(\cs[3]_net_1 ), .B(N_173), .Y(N_185));
    
endmodule


module off_on_coder_3(
       i_7,
       i_8,
       count_9,
       GLA,
       dump_state_0_off_start,
       state1ms_choice_0_reset_out
    );
output [1:1] i_7;
output [0:0] i_8;
input  [4:0] count_9;
input  GLA;
input  dump_state_0_off_start;
input  state1ms_choice_0_reset_out;

    wire \i_0_1[1] , \i_RNO_3[1] , N_17, \i_RNO_4[0] , GND, VCC, GND_0, 
        VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \i_RNO_1[1]  (.A(count_9[1]), .B(count_9[0]), .Y(N_17));
    DFN1 \i[1]  (.D(\i_RNO_3[1] ), .CLK(GLA), .Q(i_7[1]));
    GND GND_i_0 (.Y(GND_0));
    NOR3C \i_RNO[1]  (.A(\i_0_1[1] ), .B(N_17), .C(
        state1ms_choice_0_reset_out), .Y(\i_RNO_3[1] ));
    VCC VCC_i (.Y(VCC));
    NOR3B \i_RNO_0[1]  (.A(count_9[2]), .B(count_9[4]), .C(count_9[3]), 
        .Y(\i_0_1[1] ));
    NOR2B \i_RNO[0]  (.A(state1ms_choice_0_reset_out), .B(
        dump_state_0_off_start), .Y(\i_RNO_4[0] ));
    DFN1 \i[0]  (.D(\i_RNO_4[0] ), .CLK(GLA), .Q(i_8[0]));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_3(
       i_6,
       i_7,
       GLA,
       DUMP_0_dump_on,
       off_on_state_1_state_over,
       state1ms_choice_0_reset_out
    );
input  [1:1] i_6;
input  [0:0] i_7;
input  GLA;
output DUMP_0_dump_on;
output off_on_state_1_state_over;
input  state1ms_choice_0_reset_out;

    wire state_over_1_0, state_over_RNO_0_net_1, N_42, \cs_ns[1] , 
        \cs[1]_net_1 , \cs_nsss[1] , \cs_nsss[0] , GND, VCC, GND_0, 
        VCC_0;
    
    NOR2B state_over_RNO_0 (.A(i_7[0]), .B(state1ms_choice_0_reset_out)
        , .Y(state_over_1_0));
    DFN1 state_over (.D(state_over_RNO_0_net_1), .CLK(GLA), .Q(
        off_on_state_1_state_over));
    DFN1 \cs[0]  (.D(\cs_nsss[0] ), .CLK(GLA), .Q(DUMP_0_dump_on));
    NOR3C \cs_RNO[0]  (.A(N_42), .B(state1ms_choice_0_reset_out), .C(
        i_7[0]), .Y(\cs_nsss[0] ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 \cs[1]  (.D(\cs_nsss[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3C \cs_RNO[1]  (.A(\cs_ns[1] ), .B(state1ms_choice_0_reset_out), 
        .C(i_7[0]), .Y(\cs_nsss[1] ));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    MX2 \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_6[1]), .S(
        DUMP_0_dump_on), .Y(\cs_ns[1] ));
    AOI1 \cs_RNIAKJD[1]  (.A(DUMP_0_dump_on), .B(i_6[1]), .C(
        \cs[1]_net_1 ), .Y(N_42));
    AO1B state_over_RNO (.A(off_on_state_1_state_over), .B(N_42), .C(
        state_over_1_0), .Y(state_over_RNO_0_net_1));
    
endmodule


module off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_4(
       i_7,
       i_8,
       GLA,
       DUMP_0_dump_off,
       off_on_state_0_state_over,
       state1ms_choice_0_reset_out
    );
input  [1:1] i_7;
input  [0:0] i_8;
input  GLA;
output DUMP_0_dump_off;
output off_on_state_0_state_over;
input  state1ms_choice_0_reset_out;

    wire state_over_1_0, N_14, N_42, \cs_ns[1] , \cs[1]_net_1 , 
        \cs_nsss[1] , \cs_nsss[0] , GND, VCC, GND_0, VCC_0;
    
    NOR2B state_over_RNO_0 (.A(i_8[0]), .B(state1ms_choice_0_reset_out)
        , .Y(state_over_1_0));
    DFN1 state_over (.D(N_14), .CLK(GLA), .Q(off_on_state_0_state_over)
        );
    DFN1 \cs[0]  (.D(\cs_nsss[0] ), .CLK(GLA), .Q(DUMP_0_dump_off));
    NOR3C \cs_RNO[0]  (.A(N_42), .B(state1ms_choice_0_reset_out), .C(
        i_8[0]), .Y(\cs_nsss[0] ));
    AOI1 \cs_RNITUHD[1]  (.A(DUMP_0_dump_off), .B(i_7[1]), .C(
        \cs[1]_net_1 ), .Y(N_42));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 \cs[1]  (.D(\cs_nsss[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3C \cs_RNO[1]  (.A(\cs_ns[1] ), .B(state1ms_choice_0_reset_out), 
        .C(i_8[0]), .Y(\cs_nsss[1] ));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    MX2 \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_7[1]), .S(
        DUMP_0_dump_off), .Y(\cs_ns[1] ));
    AO1B state_over_RNO (.A(off_on_state_0_state_over), .B(N_42), .C(
        state_over_1_0), .Y(N_14));
    
endmodule


module dump_coder(
       i_0,
       i_1,
       i_5,
       i_8,
       i_9,
       count_3,
       dump_cho,
       dumpdata,
       count_8,
       count_1,
       GLA,
       bri_div_start_0,
       state1ms_choice_0_bri_cycle,
       top_code_0_dumpload,
       state1ms_choice_0_dump_start,
       state1ms_choice_0_reset_out
    );
output [8:6] i_0;
output [5:4] i_1;
output [3:2] i_5;
output [1:1] i_8;
output [0:0] i_9;
input  [7:5] count_3;
input  [2:0] dump_cho;
input  [11:0] dumpdata;
input  [4:0] count_8;
input  [11:8] count_1;
input  GLA;
input  bri_div_start_0;
input  state1ms_choice_0_bri_cycle;
input  top_code_0_dumpload;
input  state1ms_choice_0_dump_start;
input  state1ms_choice_0_reset_out;

    wire \i_0_0_a2_12[3] , \un1_count_3_i[0] , \i_0_0_a2_10[3] , 
        \un1_count_2_NE[0] , \i_0_0_a2_7[3] , \i_0_0_a2_6[3] , 
        \i_0_0_a2_8[3] , \i_RNO_11[3]_net_1 , \un1_count_4_5_i_0[0] , 
        \i_0_0_a2_5[3] , \i_RNO_5[3]_net_1 , \un1_count_4_0_i_0[0] , 
        \i_0_0_a2_3[3] , \un1_count_4_7_i_0[0] , 
        \un1_count_4_1_i_0[0] , \i_0_0_a2_1[3] , \para1[9]_net_1 , 
        \un1_count_4_10_i_0[0] , \para1[3]_net_1 , \i_RNO_14[3]_net_1 , 
        \para1[8]_net_1 , \un1_count_4_11_i_0[0] , \i_0_0_a2_0[4] , 
        \i_reg16_NE_8[0] , \para6_RNI7MA7[6]_net_1 , \i_reg16_5_i[0] , 
        \i_reg16_NE_5[0] , \i_reg16_NE_7[0] , \para6_RNIVL97[2]_net_1 , 
        \i_reg16_0_i[0] , \i_reg16_NE_3[0] , \i_reg16_NE_6[0] , 
        \i_reg16_7_i[0] , \i_reg16_1_i[0] , \i_reg16_NE_1[0] , 
        \para6[9]_net_1 , \i_reg16_10_i[0] , \para6[3]_net_1 , 
        \para6_RNI36A7[4]_net_1 , \para6[8]_net_1 , \i_reg16_11_i[0] , 
        \un1_count_NE_8[0] , \para5_RNI46A7[6]_net_1 , 
        \un1_count_5_i[0] , \un1_count_NE_5[0] , \un1_count_NE_7[0] , 
        \para5_RNIS597[2]_net_1 , \un1_count_0_i[0] , 
        \un1_count_NE_3[0] , \un1_count_NE_6[0] , \un1_count_7_i[0] , 
        \un1_count_1_0_i[0] , \un1_count_NE_1[0] , \para5[9]_net_1 , 
        \un1_count_10_i[0] , \para5[3]_net_1 , 
        \para5_RNI0M97[4]_net_1 , \para5[8]_net_1 , 
        \un1_count_11_i[0] , \un1_count_1_NE_8[0] , 
        \para4_RNI1M97[6]_net_1 , \un1_count_1_5_i[0] , 
        \un1_count_1_NE_5[0] , \un1_count_1_NE_7[0] , 
        \para4_RNIPL87[2]_net_1 , \un1_count_1_0_0_i[0] , 
        \un1_count_1_NE_3[0] , \un1_count_1_NE_6[0] , 
        \un1_count_1_7_i[0] , \un1_count_1_1_i[0] , 
        \un1_count_1_NE_1[0] , \para4[9]_net_1 , \un1_count_1_10_i[0] , 
        \para4[3]_net_1 , \para4_RNIT597[4]_net_1 , \para4[8]_net_1 , 
        \un1_count_1_11_i[0] , \un1_count_2_NE_8[0] , 
        \para3_RNIU597[6]_net_1 , \un1_count_2_5_i[0] , 
        \un1_count_2_NE_5[0] , \un1_count_2_NE_7[0] , 
        \para3_RNIM587[2]_net_1 , \un1_count_2_0_0_i[0] , 
        \un1_count_2_NE_3[0] , \un1_count_2_NE_6[0] , 
        \un1_count_2_7_i[0] , \un1_count_2_1_i[0] , 
        \un1_count_2_NE_1[0] , \para3[9]_net_1 , \un1_count_2_10_i[0] , 
        \para3[3]_net_1 , \para3_RNIQL87[4]_net_1 , \para3[8]_net_1 , 
        \un1_count_2_11_i[0] , \un1_count_3_NE_8[0] , 
        \para2_RNIRL87[6]_net_1 , \un1_count_3_5_i[0] , 
        \un1_count_3_NE_5[0] , \un1_count_3_NE_7[0] , 
        \para2_RNIJL77[2]_net_1 , \un1_count_3_0_0_i[0] , 
        \un1_count_3_NE_3[0] , \un1_count_3_NE_6[0] , 
        \un1_count_3_7_i[0] , \un1_count_3_1_i[0] , 
        \un1_count_3_NE_1[0] , \para2[9]_net_1 , \un1_count_3_10_i[0] , 
        \para2[3]_net_1 , \para2_RNIN587[4]_net_1 , \para2[8]_net_1 , 
        \un1_count_3_11_i[0] , \para5_4[7] , N_51, \i_RNO_3[3]_net_1 , 
        N_24, \un1_count_1_NE[0] , \i_RNO_1[4] , \un1_count_NE[0] , 
        \i_reg16_NE[0] , \para1[11]_net_1 , \para5[11]_net_1 , 
        \para4[11]_net_1 , \para3[11]_net_1 , \para2[11]_net_1 , 
        \para1[10]_net_1 , \para6[10]_net_1 , \para5[10]_net_1 , 
        \para4[10]_net_1 , \para3[10]_net_1 , \para2[10]_net_1 , 
        \para1[7]_net_1 , \para6[7]_net_1 , \para5[7]_net_1 , 
        \para4[7]_net_1 , \para3[7]_net_1 , \para2[7]_net_1 , 
        \para1[6]_net_1 , \para5[6]_net_1 , \para4[6]_net_1 , 
        \para3[6]_net_1 , \para2[6]_net_1 , \para1[5]_net_1 , 
        \para5[5]_net_1 , \para4[5]_net_1 , \para3[5]_net_1 , 
        \para2[5]_net_1 , \para1[4]_net_1 , \para5[4]_net_1 , 
        \para4[4]_net_1 , \para3[4]_net_1 , \para2[4]_net_1 , 
        \para1[2]_net_1 , \para5[2]_net_1 , \para4[2]_net_1 , 
        \para3[2]_net_1 , \para2[2]_net_1 , \para1[1]_net_1 , 
        \para5[1]_net_1 , \para4[1]_net_1 , \para3[1]_net_1 , 
        \para2[1]_net_1 , \para1[0]_net_1 , \para5[0]_net_1 , 
        \para4[0]_net_1 , \para3[0]_net_1 , \para2[0]_net_1 , 
        \i_RNO_1[5] , \i_RNO_0[6] , N_4, N_14, \para4_4[7] , 
        \para6_4[7] , \para6_4[9] , \para6_4[10] , \para6_4[11] , N_60, 
        N_59_1, N_59, N_63_1, N_280, N_61, N_12, N_53, \para6_4[3] , 
        N_8, N_6, N_57, N_58, \para6_4[8] , \para6_4[6] , \para6_4[5] , 
        \para6_4[4] , \para6_4[2] , \para6_4[1] , \para6_4[0] , 
        \para4_4[11] , \para4_4[10] , \para4_4[9] , \para4_4[8] , 
        \para4_4[6] , \para4_4[5] , \para4_4[4] , \para4_4[3] , 
        \para4_4[2] , \para4_4[1] , \para4_4[0] , \para5_4[11] , 
        \para5_4[10] , \para5_4[9] , \para5_4[3] , \i_RNO_0[8] , 
        \para6[0]_net_1 , \para6[1]_net_1 , \para6[2]_net_1 , 
        \para6[4]_net_1 , \para6[5]_net_1 , \para6[6]_net_1 , 
        \para6[11]_net_1 , GND, VCC, GND_0, VCC_0;
    
    NOR2A \i_RNO[6]  (.A(N_24), .B(\un1_count_1_NE[0] ), .Y(
        \i_RNO_0[6] ));
    NOR3C un1_para114_5_i_a2 (.A(top_code_0_dumpload), .B(dump_cho[2]), 
        .C(dump_cho[1]), .Y(N_61));
    DFN1E1 \para4[11]  (.D(\para4_4[11] ), .CLK(GLA), .E(N_59), .Q(
        \para4[11]_net_1 ));
    NOR2B \i_RNO[2]  (.A(state1ms_choice_0_reset_out), .B(
        state1ms_choice_0_bri_cycle), .Y(N_8));
    NOR2A \para4_4_0_a2[10]  (.A(dumpdata[10]), .B(dump_cho[2]), .Y(
        \para4_4[10] ));
    XNOR2 \para4_RNIND87[1]  (.A(count_8[1]), .B(\para4[1]_net_1 ), .Y(
        \un1_count_1_1_i[0] ));
    DFN1 \i[7]  (.D(N_14), .CLK(GLA), .Q(i_0[7]));
    XNOR2 \para5_RNI4VMB[10]  (.A(count_1[10]), .B(\para5[10]_net_1 ), 
        .Y(\un1_count_10_i[0] ));
    DFN1E1 \para6[1]  (.D(\para6_4[1] ), .CLK(GLA), .E(N_57), .Q(
        \para6[1]_net_1 ));
    XNOR2 \para2_RNIF577[0]  (.A(count_8[0]), .B(\para2[0]_net_1 ), .Y(
        \un1_count_3_0_0_i[0] ));
    XNOR2 \para2_RNIPD87[5]  (.A(count_3[5]), .B(\para2[5]_net_1 ), .Y(
        \un1_count_3_5_i[0] ));
    DFN1E1 \para6[7]  (.D(\para6_4[7] ), .CLK(GLA), .E(N_57), .Q(
        \para6[7]_net_1 ));
    XNOR2 \para3_RNIQL87[4]  (.A(count_8[4]), .B(\para3[4]_net_1 ), .Y(
        \para3_RNIQL87[4]_net_1 ));
    XNOR2 \para2_RNITT87[7]  (.A(count_3[7]), .B(\para2[7]_net_1 ), .Y(
        \un1_count_3_7_i[0] ));
    NOR3C \para6_RNI62O11[5]  (.A(\para6_RNI7MA7[6]_net_1 ), .B(
        \i_reg16_5_i[0] ), .C(\i_reg16_NE_5[0] ), .Y(\i_reg16_NE_8[0] )
        );
    DFN1E1 \para4[8]  (.D(\para4_4[8] ), .CLK(GLA), .E(N_59), .Q(
        \para4[8]_net_1 ));
    DFN1E1 \para2[8]  (.D(\para6_4[8] ), .CLK(GLA), .E(N_12), .Q(
        \para2[8]_net_1 ));
    XA1A \para5_RNIET1J[9]  (.A(\para5[9]_net_1 ), .B(count_1[9]), .C(
        \un1_count_10_i[0] ), .Y(\un1_count_NE_5[0] ));
    DFN1 \i[0]  (.D(N_4), .CLK(GLA), .Q(i_9[0]));
    OR3C \para4_RNI41A03[0]  (.A(\un1_count_1_NE_7[0] ), .B(
        \un1_count_1_NE_6[0] ), .C(\un1_count_1_NE_8[0] ), .Y(
        \un1_count_1_NE[0] ));
    NOR2A \para4_4_0_a2[11]  (.A(dumpdata[11]), .B(dump_cho[2]), .Y(
        \para4_4[11] ));
    XNOR2 \para6_RNIDFNB[10]  (.A(count_1[10]), .B(\para6[10]_net_1 ), 
        .Y(\i_reg16_10_i[0] ));
    NOR3C \i_RNO[3]  (.A(N_24), .B(\un1_count_1_NE[0] ), .C(
        \i_0_0_a2_12[3] ), .Y(\i_RNO_3[3]_net_1 ));
    NOR2A \para4_4_0_a2[6]  (.A(dumpdata[6]), .B(dump_cho[2]), .Y(
        \para4_4[6] ));
    NOR3C \para6_RNIUV6T[0]  (.A(\para6_RNIVL97[2]_net_1 ), .B(
        \i_reg16_0_i[0] ), .C(\i_reg16_NE_3[0] ), .Y(\i_reg16_NE_7[0] )
        );
    OA1B un1_para114_3_i_a2 (.A(dump_cho[0]), .B(dump_cho[2]), .C(
        N_59_1), .Y(N_59));
    XNOR2 \para3_RNIIL77[0]  (.A(count_8[0]), .B(\para3[0]_net_1 ), .Y(
        \un1_count_2_0_0_i[0] ));
    NOR3C \para6_RNI02N11[1]  (.A(\i_reg16_7_i[0] ), .B(
        \i_reg16_1_i[0] ), .C(\i_reg16_NE_1[0] ), .Y(\i_reg16_NE_6[0] )
        );
    NOR2A \para4_4_0_a2[9]  (.A(dumpdata[9]), .B(dump_cho[2]), .Y(
        \para4_4[9] ));
    XNOR2 \i_RNO_12[3]  (.A(count_3[5]), .B(\para1[5]_net_1 ), .Y(
        \un1_count_4_5_i_0[0] ));
    NOR3B \i_RNO[5]  (.A(N_24), .B(\un1_count_1_NE[0] ), .C(
        \un1_count_2_NE[0] ), .Y(\i_RNO_1[5] ));
    NOR3B \i_RNO[4]  (.A(N_24), .B(\un1_count_1_NE[0] ), .C(
        \i_0_0_a2_0[4] ), .Y(\i_RNO_1[4] ));
    NOR3C \i_RNO_1[3]  (.A(\i_0_0_a2_7[3] ), .B(\i_0_0_a2_6[3] ), .C(
        \i_0_0_a2_8[3] ), .Y(\i_0_0_a2_10[3] ));
    XNOR2 \para3_RNIKT77[1]  (.A(count_8[1]), .B(\para3[1]_net_1 ), .Y(
        \un1_count_2_1_i[0] ));
    DFN1E1 \para2[10]  (.D(\para6_4[10] ), .CLK(GLA), .E(N_12), .Q(
        \para2[10]_net_1 ));
    OR3C \para6_RNI44M03[0]  (.A(\i_reg16_NE_7[0] ), .B(
        \i_reg16_NE_6[0] ), .C(\i_reg16_NE_8[0] ), .Y(\i_reg16_NE[0] ));
    NOR2A \para2_4_0_a2[7]  (.A(dumpdata[7]), .B(dump_cho[1]), .Y(
        \para6_4[7] ));
    DFN1E1 \para1[9]  (.D(\para4_4[9] ), .CLK(GLA), .E(N_280), .Q(
        \para1[9]_net_1 ));
    XNOR2 \para3_RNIM587[2]  (.A(count_8[2]), .B(\para3[2]_net_1 ), .Y(
        \para3_RNIM587[2]_net_1 ));
    DFN1E1 \para1[8]  (.D(\para4_4[8] ), .CLK(GLA), .E(N_280), .Q(
        \para1[8]_net_1 ));
    XA1A \para6_RNIQT2J[9]  (.A(\para6[9]_net_1 ), .B(count_1[9]), .C(
        \i_reg16_10_i[0] ), .Y(\i_reg16_NE_5[0] ));
    DFN1E1 \para5[5]  (.D(\para6_4[5] ), .CLK(GLA), .E(N_58), .Q(
        \para5[5]_net_1 ));
    NOR3C \para3_RNIA0H11[1]  (.A(\un1_count_2_7_i[0] ), .B(
        \un1_count_2_1_i[0] ), .C(\un1_count_2_NE_1[0] ), .Y(
        \un1_count_2_NE_6[0] ));
    DFN1E1 \para4[10]  (.D(\para4_4[10] ), .CLK(GLA), .E(N_59), .Q(
        \para4[10]_net_1 ));
    NOR3C \para5_RNIK1M11[5]  (.A(\para5_RNI46A7[6]_net_1 ), .B(
        \un1_count_5_i[0] ), .C(\un1_count_NE_5[0] ), .Y(
        \un1_count_NE_8[0] ));
    DFN1E1 \para3[3]  (.D(\para4_4[3] ), .CLK(GLA), .E(N_60), .Q(
        \para3[3]_net_1 ));
    DFN1E1 \para6[0]  (.D(\para6_4[0] ), .CLK(GLA), .E(N_57), .Q(
        \para6[0]_net_1 ));
    XA1A \i_RNO_13[3]  (.A(\para1[9]_net_1 ), .B(count_1[9]), .C(
        \un1_count_4_10_i_0[0] ), .Y(\i_0_0_a2_5[3] ));
    NOR2A un1_para114_6_i_a2_1 (.A(top_code_0_dumpload), .B(
        dump_cho[2]), .Y(N_63_1));
    XA1A \para6_RNI44KE[3]  (.A(\para6[3]_net_1 ), .B(count_8[3]), .C(
        \para6_RNI36A7[4]_net_1 ), .Y(\i_reg16_NE_3[0] ));
    DFN1E1 \para3[7]  (.D(\para4_4[7] ), .CLK(GLA), .E(N_60), .Q(
        \para3[7]_net_1 ));
    XA1A \para3_RNIMKVI[8]  (.A(\para3[8]_net_1 ), .B(count_1[8]), .C(
        \un1_count_2_11_i[0] ), .Y(\un1_count_2_NE_1[0] ));
    NOR2A \para2_4_0_a2[2]  (.A(dumpdata[2]), .B(dump_cho[1]), .Y(
        \para6_4[2] ));
    NOR2B \i_RNO[0]  (.A(state1ms_choice_0_reset_out), .B(
        state1ms_choice_0_dump_start), .Y(N_4));
    NOR2A \para4_4_0_a2[8]  (.A(dumpdata[8]), .B(dump_cho[2]), .Y(
        \para4_4[8] ));
    XNOR2 \para2_RNIBELB[11]  (.A(count_1[11]), .B(\para2[11]_net_1 ), 
        .Y(\un1_count_3_11_i[0] ));
    XNOR2 \i_RNO_16[3]  (.A(count_1[10]), .B(\para1[10]_net_1 ), .Y(
        \un1_count_4_10_i_0[0] ));
    NOR2 un1_para114_i_o2 (.A(dump_cho[1]), .B(dump_cho[0]), .Y(N_51));
    XNOR2 \para5_RNIS597[2]  (.A(count_8[2]), .B(\para5[2]_net_1 ), .Y(
        \para5_RNIS597[2]_net_1 ));
    NOR2A \para2_4_0_a2[5]  (.A(dumpdata[5]), .B(dump_cho[1]), .Y(
        \para6_4[5] ));
    GND GND_i (.Y(GND));
    XA1A \i_RNO_10[3]  (.A(\para1[8]_net_1 ), .B(count_1[8]), .C(
        \un1_count_4_11_i_0[0] ), .Y(\i_0_0_a2_1[3] ));
    DFN1E1 \para3[11]  (.D(\para4_4[11] ), .CLK(GLA), .E(N_60), .Q(
        \para3[11]_net_1 ));
    DFN1E1 \para2[9]  (.D(\para6_4[9] ), .CLK(GLA), .E(N_12), .Q(
        \para2[9]_net_1 ));
    NOR3C \para5_RNIIV4T[0]  (.A(\para5_RNIS597[2]_net_1 ), .B(
        \un1_count_0_i[0] ), .C(\un1_count_NE_3[0] ), .Y(
        \un1_count_NE_7[0] ));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR3C \para2_RNIOVE11[1]  (.A(\un1_count_3_7_i[0] ), .B(
        \un1_count_3_1_i[0] ), .C(\un1_count_3_NE_1[0] ), .Y(
        \un1_count_3_NE_6[0] ));
    XNOR2 \para3_RNIU597[6]  (.A(count_3[6]), .B(\para3[6]_net_1 ), .Y(
        \para3_RNIU597[6]_net_1 ));
    XNOR2 \para5_RNI6VMB[11]  (.A(count_1[11]), .B(\para5[11]_net_1 ), 
        .Y(\un1_count_11_i[0] ));
    NOR2A \para4_4_0_a2[4]  (.A(dumpdata[4]), .B(dump_cho[2]), .Y(
        \para4_4[4] ));
    XNOR2 \para3_RNIST87[5]  (.A(count_3[5]), .B(\para3[5]_net_1 ), .Y(
        \un1_count_2_5_i[0] ));
    XNOR2 \i_RNO_6[3]  (.A(count_8[0]), .B(\para1[0]_net_1 ), .Y(
        \un1_count_4_0_i_0[0] ));
    NOR2B \i_RNO[1]  (.A(state1ms_choice_0_reset_out), .B(
        bri_div_start_0), .Y(N_6));
    XA1A \i_RNO_7[3]  (.A(\para1[3]_net_1 ), .B(count_8[3]), .C(
        \i_RNO_14[3]_net_1 ), .Y(\i_0_0_a2_3[3] ));
    XNOR2 \para5_RNI2U97[5]  (.A(count_3[5]), .B(\para5[5]_net_1 ), .Y(
        \un1_count_5_i[0] ));
    XNOR2 \i_RNO_14[3]  (.A(count_8[4]), .B(\para1[4]_net_1 ), .Y(
        \i_RNO_14[3]_net_1 ));
    XA1A \para4_RNI2L0J[8]  (.A(\para4[8]_net_1 ), .B(count_1[8]), .C(
        \un1_count_1_11_i[0] ), .Y(\un1_count_1_NE_1[0] ));
    XNOR2 \para4_RNITEMB[11]  (.A(count_1[11]), .B(\para4[11]_net_1 ), 
        .Y(\un1_count_1_11_i[0] ));
    XNOR2 \para3_RNIIULB[10]  (.A(count_1[10]), .B(\para3[10]_net_1 ), 
        .Y(\un1_count_2_10_i[0] ));
    DFN1E1 \para3[1]  (.D(\para4_4[1] ), .CLK(GLA), .E(N_60), .Q(
        \para3[1]_net_1 ));
    XNOR2 \para6_RNIVL97[2]  (.A(count_8[2]), .B(\para6[2]_net_1 ), .Y(
        \para6_RNIVL97[2]_net_1 ));
    DFN1E1 \para1[4]  (.D(\para4_4[4] ), .CLK(GLA), .E(N_280), .Q(
        \para1[4]_net_1 ));
    NOR3B un1_para114_i_a2 (.A(top_code_0_dumpload), .B(dump_cho[2]), 
        .C(N_51), .Y(N_57));
    XNOR2 \para2_RNI9ELB[10]  (.A(count_1[10]), .B(\para2[10]_net_1 ), 
        .Y(\un1_count_3_10_i[0] ));
    NOR2A \para2_4_0_a2[0]  (.A(dumpdata[0]), .B(dump_cho[1]), .Y(
        \para6_4[0] ));
    NOR2A un1_para114_2_i_o2 (.A(dump_cho[0]), .B(dump_cho[1]), .Y(
        N_53));
    DFN1E1 \para6[2]  (.D(\para6_4[2] ), .CLK(GLA), .E(N_57), .Q(
        \para6[2]_net_1 ));
    XNOR2 \para5_RNI6EA7[7]  (.A(count_3[7]), .B(\para5[7]_net_1 ), .Y(
        \un1_count_7_i[0] ));
    XA1A \para3_RNII3HE[3]  (.A(\para3[3]_net_1 ), .B(count_8[3]), .C(
        \para3_RNIQL87[4]_net_1 ), .Y(\un1_count_2_NE_3[0] ));
    XA1A \para4_RNI2T0J[9]  (.A(\para4[9]_net_1 ), .B(count_1[9]), .C(
        \un1_count_1_10_i[0] ), .Y(\un1_count_1_NE_5[0] ));
    XA1A \para6_RNIQL2J[8]  (.A(\para6[8]_net_1 ), .B(count_1[8]), .C(
        \i_reg16_11_i[0] ), .Y(\i_reg16_NE_1[0] ));
    DFN1E1 \para4[5]  (.D(\para4_4[5] ), .CLK(GLA), .E(N_59), .Q(
        \para4[5]_net_1 ));
    NOR2A \para4_4_0_a2[3]  (.A(dumpdata[3]), .B(dump_cho[2]), .Y(
        \para4_4[3] ));
    VCC VCC_i (.Y(VCC));
    DFN1E1 \para2[6]  (.D(\para6_4[6] ), .CLK(GLA), .E(N_12), .Q(
        \para2[6]_net_1 ));
    XNOR2 \para3_RNI0E97[7]  (.A(count_3[7]), .B(\para3[7]_net_1 ), .Y(
        \un1_count_2_7_i[0] ));
    DFN1E1 \para2[3]  (.D(\para6_4[3] ), .CLK(GLA), .E(N_12), .Q(
        \para2[3]_net_1 ));
    DFN1E1 \para2[5]  (.D(\para6_4[5] ), .CLK(GLA), .E(N_12), .Q(
        \para2[5]_net_1 ));
    NOR2A \para4_4_0_a2[1]  (.A(dumpdata[1]), .B(dump_cho[2]), .Y(
        \para4_4[1] ));
    DFN1E1 \para3[8]  (.D(\para4_4[8] ), .CLK(GLA), .E(N_60), .Q(
        \para3[8]_net_1 ));
    XNOR2 \para6_RNI7MA7[6]  (.A(count_3[6]), .B(\para6[6]_net_1 ), .Y(
        \para6_RNI7MA7[6]_net_1 ));
    XNOR2 \para4_RNIT597[4]  (.A(count_8[4]), .B(\para4[4]_net_1 ), .Y(
        \para4_RNIT597[4]_net_1 ));
    DFN1E1 \para6[6]  (.D(\para6_4[6] ), .CLK(GLA), .E(N_57), .Q(
        \para6[6]_net_1 ));
    XNOR2 \para5_RNIQT87[1]  (.A(count_8[1]), .B(\para5[1]_net_1 ), .Y(
        \un1_count_1_0_i[0] ));
    DFN1E1 \para4[0]  (.D(\para4_4[0] ), .CLK(GLA), .E(N_59), .Q(
        \para4[0]_net_1 ));
    OR3C \para5_RNIK2G03[0]  (.A(\un1_count_NE_7[0] ), .B(
        \un1_count_NE_6[0] ), .C(\un1_count_NE_8[0] ), .Y(
        \un1_count_NE[0] ));
    DFN1E1 \para3[10]  (.D(\para4_4[10] ), .CLK(GLA), .E(N_60), .Q(
        \para3[10]_net_1 ));
    DFN1E1 \para6[9]  (.D(\para6_4[9] ), .CLK(GLA), .E(N_57), .Q(
        \para6[9]_net_1 ));
    DFN1E1 \para5[8]  (.D(\para6_4[8] ), .CLK(GLA), .E(N_58), .Q(
        \para5[8]_net_1 ));
    DFN1E1 \para1[3]  (.D(\para4_4[3] ), .CLK(GLA), .E(N_280), .Q(
        \para1[3]_net_1 ));
    DFN1E1 \para1[2]  (.D(\para4_4[2] ), .CLK(GLA), .E(N_280), .Q(
        \para1[2]_net_1 ));
    DFN1E1 \para3[6]  (.D(\para4_4[6] ), .CLK(GLA), .E(N_60), .Q(
        \para3[6]_net_1 ));
    OR2B un1_para114_4_i_a2_1 (.A(dump_cho[1]), .B(top_code_0_dumpload)
        , .Y(N_59_1));
    XA1A \para4_RNIO3IE[3]  (.A(\para4[3]_net_1 ), .B(count_8[3]), .C(
        \para4_RNIT597[4]_net_1 ), .Y(\un1_count_1_NE_3[0] ));
    DFN1E1 \para4[2]  (.D(\para4_4[2] ), .CLK(GLA), .E(N_59), .Q(
        \para4[2]_net_1 ));
    NOR3C \para3_RNIQU0T[0]  (.A(\para3_RNIM587[2]_net_1 ), .B(
        \un1_count_2_0_0_i[0] ), .C(\un1_count_2_NE_3[0] ), .Y(
        \un1_count_2_NE_7[0] ));
    XNOR2 \para4_RNIVD97[5]  (.A(count_3[5]), .B(\para4[5]_net_1 ), .Y(
        \un1_count_1_5_i[0] ));
    DFN1E1 \para2[4]  (.D(\para6_4[4] ), .CLK(GLA), .E(N_12), .Q(
        \para2[4]_net_1 ));
    XA1A \para2_RNIAKUI[8]  (.A(\para2[8]_net_1 ), .B(count_1[8]), .C(
        \un1_count_3_11_i[0] ), .Y(\un1_count_3_NE_1[0] ));
    DFN1E1 \para1[11]  (.D(\para4_4[11] ), .CLK(GLA), .E(N_280), .Q(
        \para1[11]_net_1 ));
    DFN1E1 \para6[4]  (.D(\para6_4[4] ), .CLK(GLA), .E(N_57), .Q(
        \para6[4]_net_1 ));
    DFN1E1 \para5[11]  (.D(\para5_4[11] ), .CLK(GLA), .E(N_58), .Q(
        \para5[11]_net_1 ));
    XNOR2 \para5_RNIOL87[0]  (.A(count_8[0]), .B(\para5[0]_net_1 ), .Y(
        \un1_count_0_i[0] ));
    DFN1E1 \para5[4]  (.D(\para6_4[4] ), .CLK(GLA), .E(N_58), .Q(
        \para5[4]_net_1 ));
    NOR3C \para4_RNI6V2T[0]  (.A(\para4_RNIPL87[2]_net_1 ), .B(
        \un1_count_1_0_0_i[0] ), .C(\un1_count_1_NE_3[0] ), .Y(
        \un1_count_1_NE_7[0] ));
    DFN1E1 \para4[3]  (.D(\para4_4[3] ), .CLK(GLA), .E(N_59), .Q(
        \para4[3]_net_1 ));
    NOR3C \para3_RNIG0I11[5]  (.A(\para3_RNIU597[6]_net_1 ), .B(
        \un1_count_2_5_i[0] ), .C(\un1_count_2_NE_5[0] ), .Y(
        \un1_count_2_NE_8[0] ));
    XA1A \para5_RNIU3JE[3]  (.A(\para5[3]_net_1 ), .B(count_8[3]), .C(
        \para5_RNI0M97[4]_net_1 ), .Y(\un1_count_NE_3[0] ));
    DFN1E1 \para6[11]  (.D(\para6_4[11] ), .CLK(GLA), .E(N_57), .Q(
        \para6[11]_net_1 ));
    XNOR2 \para2_RNIRL87[6]  (.A(count_3[6]), .B(\para2[6]_net_1 ), .Y(
        \para2_RNIRL87[6]_net_1 ));
    DFN1E1 \para6[5]  (.D(\para6_4[5] ), .CLK(GLA), .E(N_57), .Q(
        \para6[5]_net_1 ));
    DFN1E1 \para3[4]  (.D(\para4_4[4] ), .CLK(GLA), .E(N_60), .Q(
        \para3[4]_net_1 ));
    DFN1 \i[2]  (.D(N_8), .CLK(GLA), .Q(i_5[2]));
    DFN1E1 \para1[6]  (.D(\para4_4[6] ), .CLK(GLA), .E(N_280), .Q(
        \para1[6]_net_1 ));
    XNOR2 \i_RNO_5[3]  (.A(count_8[2]), .B(\para1[2]_net_1 ), .Y(
        \i_RNO_5[3]_net_1 ));
    DFN1E1 \para4[4]  (.D(\para4_4[4] ), .CLK(GLA), .E(N_59), .Q(
        \para4[4]_net_1 ));
    OR3C \para3_RNIKV303[0]  (.A(\un1_count_2_NE_7[0] ), .B(
        \un1_count_2_NE_6[0] ), .C(\un1_count_2_NE_8[0] ), .Y(
        \un1_count_2_NE[0] ));
    XNOR2 \para6_RNI5EA7[5]  (.A(count_3[5]), .B(\para6[5]_net_1 ), .Y(
        \i_reg16_5_i[0] ));
    DFN1E1 \para1[5]  (.D(\para4_4[5] ), .CLK(GLA), .E(N_280), .Q(
        \para1[5]_net_1 ));
    DFN1E1 \para5[3]  (.D(\para5_4[3] ), .CLK(GLA), .E(N_58), .Q(
        \para5[3]_net_1 ));
    DFN1E1 \para2[7]  (.D(\para6_4[7] ), .CLK(GLA), .E(N_12), .Q(
        \para2[7]_net_1 ));
    NOR2A \para2_4_0_a2[6]  (.A(dumpdata[6]), .B(dump_cho[1]), .Y(
        \para6_4[6] ));
    OA1C un1_para114_4_i_a2 (.A(dump_cho[0]), .B(dump_cho[2]), .C(
        N_59_1), .Y(N_60));
    DFN1E1 \para4[7]  (.D(\para4_4[7] ), .CLK(GLA), .E(N_59), .Q(
        \para4[7]_net_1 ));
    XA1A \para2_RNIASUI[9]  (.A(\para2[9]_net_1 ), .B(count_1[9]), .C(
        \un1_count_3_10_i[0] ), .Y(\un1_count_3_NE_5[0] ));
    XNOR2 \i_RNO_8[3]  (.A(count_3[7]), .B(\para1[7]_net_1 ), .Y(
        \un1_count_4_7_i_0[0] ));
    XNOR2 \para2_RNIJL77[2]  (.A(count_8[2]), .B(\para2[2]_net_1 ), .Y(
        \para2_RNIJL77[2]_net_1 ));
    XNOR2 \para4_RNI1M97[6]  (.A(count_3[6]), .B(\para4[6]_net_1 ), .Y(
        \para4_RNI1M97[6]_net_1 ));
    NOR2A \para2_4_0_a2[9]  (.A(dumpdata[9]), .B(dump_cho[1]), .Y(
        \para6_4[9] ));
    AO1 un1_para114_6_i (.A(N_63_1), .B(N_51), .C(N_61), .Y(N_280));
    XNOR2 \para5_RNI0M97[4]  (.A(count_8[4]), .B(\para5[4]_net_1 ), .Y(
        \para5_RNI0M97[4]_net_1 ));
    DFN1 \i[6]  (.D(\i_RNO_0[6] ), .CLK(GLA), .Q(i_0[6]));
    XNOR2 \i_RNO_11[3]  (.A(count_3[6]), .B(\para1[6]_net_1 ), .Y(
        \i_RNO_11[3]_net_1 ));
    DFN1E1 \para2[0]  (.D(\para6_4[0] ), .CLK(GLA), .E(N_12), .Q(
        \para2[0]_net_1 ));
    DFN1 \i[4]  (.D(\i_RNO_1[4] ), .CLK(GLA), .Q(i_1[4]));
    DFN1E1 \para5[0]  (.D(\para6_4[0] ), .CLK(GLA), .E(N_58), .Q(
        \para5[0]_net_1 ));
    DFN1E1 \para5[2]  (.D(\para6_4[2] ), .CLK(GLA), .E(N_58), .Q(
        \para5[2]_net_1 ));
    NOR2A \para4_4_0_a2[7]  (.A(dumpdata[7]), .B(dump_cho[2]), .Y(
        \para4_4[7] ));
    NOR2B \para5_RNO[10]  (.A(dumpdata[10]), .B(N_51), .Y(
        \para5_4[10] ));
    GND GND_i_0 (.Y(GND_0));
    DFN1E1 \para1[0]  (.D(\para4_4[0] ), .CLK(GLA), .E(N_280), .Q(
        \para1[0]_net_1 ));
    XNOR2 \para4_RNIL587[0]  (.A(count_8[0]), .B(\para4[0]_net_1 ), .Y(
        \un1_count_1_0_0_i[0] ));
    NOR3C \para2_RNIEUUS[0]  (.A(\para2_RNIJL77[2]_net_1 ), .B(
        \un1_count_3_0_0_i[0] ), .C(\un1_count_3_NE_3[0] ), .Y(
        \un1_count_3_NE_7[0] ));
    DFN1E1 \para1[10]  (.D(\para4_4[10] ), .CLK(GLA), .E(N_280), .Q(
        \para1[10]_net_1 ));
    XNOR2 \para4_RNI3U97[7]  (.A(count_3[7]), .B(\para4[7]_net_1 ), .Y(
        \un1_count_1_7_i[0] ));
    DFN1E1 \para5[10]  (.D(\para5_4[10] ), .CLK(GLA), .E(N_58), .Q(
        \para5[10]_net_1 ));
    NOR3C \para4_RNIS0J11[1]  (.A(\un1_count_1_7_i[0] ), .B(
        \un1_count_1_1_i[0] ), .C(\un1_count_1_NE_1[0] ), .Y(
        \un1_count_1_NE_6[0] ));
    DFN1E1 \para1[1]  (.D(\para4_4[1] ), .CLK(GLA), .E(N_280), .Q(
        \para1[1]_net_1 ));
    NOR3B un1_para114_2_i_a2 (.A(top_code_0_dumpload), .B(dump_cho[2]), 
        .C(N_53), .Y(N_58));
    NOR3C \para5_RNO[7]  (.A(dumpdata[7]), .B(dump_cho[2]), .C(N_51), 
        .Y(\para5_4[7] ));
    DFN1E1 \para3[5]  (.D(\para4_4[5] ), .CLK(GLA), .E(N_60), .Q(
        \para3[5]_net_1 ));
    XNOR2 \para5_RNI46A7[6]  (.A(count_3[6]), .B(\para5[6]_net_1 ), .Y(
        \para5_RNI46A7[6]_net_1 ));
    DFN1E1 \para5[1]  (.D(\para6_4[1] ), .CLK(GLA), .E(N_58), .Q(
        \para5[1]_net_1 ));
    DFN1E1 \para2[2]  (.D(\para6_4[2] ), .CLK(GLA), .E(N_12), .Q(
        \para2[2]_net_1 ));
    DFN1E1 \para6[8]  (.D(\para6_4[8] ), .CLK(GLA), .E(N_57), .Q(
        \para6[8]_net_1 ));
    DFN1E1 \para6[10]  (.D(\para6_4[10] ), .CLK(GLA), .E(N_57), .Q(
        \para6[10]_net_1 ));
    XNOR2 \para6_RNI9UA7[7]  (.A(count_3[7]), .B(\para6[7]_net_1 ), .Y(
        \i_reg16_7_i[0] ));
    NOR3C \para5_RNIE1L11[1]  (.A(\un1_count_7_i[0] ), .B(
        \un1_count_1_0_i[0] ), .C(\un1_count_NE_1[0] ), .Y(
        \un1_count_NE_6[0] ));
    NOR2B \para5_RNO[3]  (.A(dumpdata[3]), .B(N_51), .Y(\para5_4[3] ));
    NOR2A \para2_4_0_a2[8]  (.A(dumpdata[8]), .B(dump_cho[1]), .Y(
        \para6_4[8] ));
    NOR2A \para4_4_0_a2[2]  (.A(dumpdata[2]), .B(dump_cho[2]), .Y(
        \para4_4[2] ));
    OR3C \para2_RNI4UTV2[0]  (.A(\un1_count_3_NE_7[0] ), .B(
        \un1_count_3_NE_6[0] ), .C(\un1_count_3_NE_8[0] ), .Y(
        \un1_count_3_i[0] ));
    NOR2A \i_RNO[8]  (.A(state1ms_choice_0_reset_out), .B(
        \i_reg16_NE[0] ), .Y(\i_RNO_0[8] ));
    DFN1E1 \para6[3]  (.D(\para6_4[3] ), .CLK(GLA), .E(N_57), .Q(
        \para6[3]_net_1 ));
    XNOR2 \para6_RNIR597[0]  (.A(count_8[0]), .B(\para6[0]_net_1 ), .Y(
        \i_reg16_0_i[0] ));
    DFN1E1 \para5[6]  (.D(\para6_4[6] ), .CLK(GLA), .E(N_58), .Q(
        \para5[6]_net_1 ));
    NOR2A \para4_4_0_a2[5]  (.A(dumpdata[5]), .B(dump_cho[2]), .Y(
        \para4_4[5] ));
    DFN1E1 \para5[7]  (.D(\para5_4[7] ), .CLK(GLA), .E(N_58), .Q(
        \para5[7]_net_1 ));
    DFN1E1 \para4[9]  (.D(\para4_4[9] ), .CLK(GLA), .E(N_59), .Q(
        \para4[9]_net_1 ));
    DFN1E1 \para3[0]  (.D(\para4_4[0] ), .CLK(GLA), .E(N_60), .Q(
        \para3[0]_net_1 ));
    NOR2A \para2_4_0_a2[4]  (.A(dumpdata[4]), .B(dump_cho[1]), .Y(
        \para6_4[4] ));
    XA1A \para3_RNIMSVI[9]  (.A(\para3[9]_net_1 ), .B(count_1[9]), .C(
        \un1_count_2_10_i[0] ), .Y(\un1_count_2_NE_5[0] ));
    NOR3C \i_RNO_4[3]  (.A(\i_RNO_11[3]_net_1 ), .B(
        \un1_count_4_5_i_0[0] ), .C(\i_0_0_a2_5[3] ), .Y(
        \i_0_0_a2_8[3] ));
    XNOR2 \para4_RNIPL87[2]  (.A(count_8[2]), .B(\para4[2]_net_1 ), .Y(
        \para4_RNIPL87[2]_net_1 ));
    DFN1 \i[5]  (.D(\i_RNO_1[5] ), .CLK(GLA), .Q(i_1[5]));
    DFN1 \i[8]  (.D(\i_RNO_0[8] ), .CLK(GLA), .Q(i_0[8]));
    DFN1E1 \para2[1]  (.D(\para6_4[1] ), .CLK(GLA), .E(N_12), .Q(
        \para2[1]_net_1 ));
    DFN1E1 \para3[2]  (.D(\para4_4[2] ), .CLK(GLA), .E(N_60), .Q(
        \para3[2]_net_1 ));
    NOR3C \para4_RNI21K11[5]  (.A(\para4_RNI1M97[6]_net_1 ), .B(
        \un1_count_1_5_i[0] ), .C(\un1_count_1_NE_5[0] ), .Y(
        \un1_count_1_NE_8[0] ));
    DFN1E1 \para4[1]  (.D(\para4_4[1] ), .CLK(GLA), .E(N_59), .Q(
        \para4[1]_net_1 ));
    XNOR2 \para3_RNIKULB[11]  (.A(count_1[11]), .B(\para3[11]_net_1 ), 
        .Y(\un1_count_2_11_i[0] ));
    XA1A \para2_RNIC3GE[3]  (.A(\para2[3]_net_1 ), .B(count_8[3]), .C(
        \para2_RNIN587[4]_net_1 ), .Y(\un1_count_3_NE_3[0] ));
    XNOR2 \para6_RNIFFNB[11]  (.A(count_1[11]), .B(\para6[11]_net_1 ), 
        .Y(\i_reg16_11_i[0] ));
    XNOR2 \para4_RNIREMB[10]  (.A(count_1[10]), .B(\para4[10]_net_1 ), 
        .Y(\un1_count_1_10_i[0] ));
    DFN1E1 \para3[9]  (.D(\para4_4[9] ), .CLK(GLA), .E(N_60), .Q(
        \para3[9]_net_1 ));
    NOR2A \para4_4_0_a2[0]  (.A(dumpdata[0]), .B(dump_cho[2]), .Y(
        \para4_4[0] ));
    OR2A \i_RNO_0[4]  (.A(\un1_count_2_NE[0] ), .B(\un1_count_3_i[0] ), 
        .Y(\i_0_0_a2_0[4] ));
    XNOR2 \para2_RNIN587[4]  (.A(count_8[4]), .B(\para2[4]_net_1 ), .Y(
        \para2_RNIN587[4]_net_1 ));
    AO1 un1_para114_5_i (.A(N_63_1), .B(N_53), .C(N_61), .Y(N_12));
    NOR2A \para2_4_0_a2[3]  (.A(dumpdata[3]), .B(dump_cho[1]), .Y(
        \para6_4[3] ));
    DFN1 \i[3]  (.D(\i_RNO_3[3]_net_1 ), .CLK(GLA), .Q(i_5[3]));
    NOR3C \i_RNO_3[3]  (.A(\un1_count_4_7_i_0[0] ), .B(
        \un1_count_4_1_i_0[0] ), .C(\i_0_0_a2_1[3] ), .Y(
        \i_0_0_a2_6[3] ));
    XA1A \para5_RNIEL1J[8]  (.A(\para5[8]_net_1 ), .B(count_1[8]), .C(
        \un1_count_11_i[0] ), .Y(\un1_count_NE_1[0] ));
    XNOR2 \para2_RNIHD77[1]  (.A(count_8[1]), .B(\para2[1]_net_1 ), .Y(
        \un1_count_3_1_i[0] ));
    NOR2A \para2_4_0_a2[1]  (.A(dumpdata[1]), .B(dump_cho[1]), .Y(
        \para6_4[1] ));
    XNOR2 \i_RNO_9[3]  (.A(count_8[1]), .B(\para1[1]_net_1 ), .Y(
        \un1_count_4_1_i_0[0] ));
    NOR2A \para2_4_0_a2[11]  (.A(dumpdata[11]), .B(dump_cho[1]), .Y(
        \para6_4[11] ));
    DFN1E1 \para4[6]  (.D(\para4_4[6] ), .CLK(GLA), .E(N_59), .Q(
        \para4[6]_net_1 ));
    NOR3C \i_RNO_0[3]  (.A(\un1_count_3_i[0] ), .B(\i_0_0_a2_10[3] ), 
        .C(\un1_count_2_NE[0] ), .Y(\i_0_0_a2_12[3] ));
    NOR2B \para5_RNO[11]  (.A(dumpdata[11]), .B(N_51), .Y(
        \para5_4[11] ));
    DFN1 \i[1]  (.D(N_6), .CLK(GLA), .Q(i_8[1]));
    NOR3B \i_RNO[7]  (.A(\i_reg16_NE[0] ), .B(
        state1ms_choice_0_reset_out), .C(\un1_count_NE[0] ), .Y(N_14));
    NOR3C \para2_RNIUVF11[5]  (.A(\para2_RNIRL87[6]_net_1 ), .B(
        \un1_count_3_5_i[0] ), .C(\un1_count_3_NE_5[0] ), .Y(
        \un1_count_3_NE_8[0] ));
    NOR2B \para5_RNO[9]  (.A(dumpdata[9]), .B(N_51), .Y(\para5_4[9] ));
    DFN1E1 \para5[9]  (.D(\para5_4[9] ), .CLK(GLA), .E(N_58), .Q(
        \para5[9]_net_1 ));
    XNOR2 \para6_RNITD97[1]  (.A(count_8[1]), .B(\para6[1]_net_1 ), .Y(
        \i_reg16_1_i[0] ));
    DFN1E1 \para2[11]  (.D(\para6_4[11] ), .CLK(GLA), .E(N_12), .Q(
        \para2[11]_net_1 ));
    DFN1E1 \para1[7]  (.D(\para4_4[7] ), .CLK(GLA), .E(N_280), .Q(
        \para1[7]_net_1 ));
    NOR3C \i_RNO_2[3]  (.A(\i_RNO_5[3]_net_1 ), .B(
        \un1_count_4_0_i_0[0] ), .C(\i_0_0_a2_3[3] ), .Y(
        \i_0_0_a2_7[3] ));
    NOR2A \para2_4_0_a2[10]  (.A(dumpdata[10]), .B(dump_cho[1]), .Y(
        \para6_4[10] ));
    XNOR2 \para6_RNI36A7[4]  (.A(count_8[4]), .B(\para6[4]_net_1 ), .Y(
        \para6_RNI36A7[4]_net_1 ));
    NOR3C \para5_RNIN5736[0]  (.A(\i_reg16_NE[0] ), .B(
        state1ms_choice_0_reset_out), .C(\un1_count_NE[0] ), .Y(N_24));
    XNOR2 \i_RNO_15[3]  (.A(count_1[11]), .B(\para1[11]_net_1 ), .Y(
        \un1_count_4_11_i_0[0] ));
    
endmodule


module dump_timer(
       count_1,
       count_8,
       count_3,
       GLA,
       state1ms_choice_0_reset_out,
       dump_state_0_timer_start,
       state1ms_choice_0_dump_start
    );
output [11:8] count_1;
output [4:0] count_8;
output [7:5] count_3;
input  GLA;
input  state1ms_choice_0_reset_out;
input  dump_state_0_timer_start;
input  state1ms_choice_0_dump_start;

    wire count_n7_0_i_0, count_0_sqmuxa_net_1, 
        \count_RNI4LSV[1]_net_1 , count_n7_0_i_o3_m3_0_a2_4, 
        count_n7_0_i_o3_m3_0_a2_1, count_n7_0_i_o3_m3_0_a2_0, 
        count_n7_0_i_o3_m3_0_a2_2, N_5, N_7, N_23, N_9, N_24, N_11, 
        N_25, N_13, N_26, N_15, N_61, N_28, N_17, N_19, count_n0, 
        count_n9, N_30, count_n10, N_31, count_n11, N_32, GND, VCC, 
        GND_0, VCC_0;
    
    DFN1 \count[5]  (.D(N_13), .CLK(GLA), .Q(count_3[5]));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_8[1]));
    DFN1 \count[10]  (.D(count_n10), .CLK(GLA), .Q(count_1[10]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_8[0]));
    AOI1 \count_RNO_0[6]  (.A(count_3[5]), .B(N_26), .C(count_3[6]), 
        .Y(N_61));
    NOR2A \count_RNIMPTB[2]  (.A(count_8[2]), .B(N_23), .Y(N_24));
    OA1B \count_RNO[7]  (.A(N_28), .B(count_3[7]), .C(count_n7_0_i_0), 
        .Y(N_17));
    NOR3C \count_RNI18UN[3]  (.A(count_n7_0_i_o3_m3_0_a2_1), .B(
        count_n7_0_i_o3_m3_0_a2_0), .C(count_n7_0_i_o3_m3_0_a2_2), .Y(
        count_n7_0_i_o3_m3_0_a2_4));
    XA1C \count_RNO[2]  (.A(N_23), .B(count_8[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR2B \count_RNIAATF[3]  (.A(count_8[3]), .B(N_24), .Y(N_25));
    XA1C \count_RNO[9]  (.A(count_1[9]), .B(N_30), .C(
        count_0_sqmuxa_net_1), .Y(count_n9));
    VCC VCC_i (.Y(VCC));
    XA1C \count_RNO[4]  (.A(N_25), .B(count_8[4]), .C(
        count_0_sqmuxa_net_1), .Y(N_11));
    DFN1 \count[8]  (.D(N_19), .CLK(GLA), .Q(count_1[8]));
    OR2A \count_RNIN2T71[9]  (.A(count_1[9]), .B(N_30), .Y(N_31));
    XA1C \count_RNO[10]  (.A(count_1[10]), .B(N_31), .C(
        count_0_sqmuxa_net_1), .Y(count_n10));
    NOR2A \count_RNIVUSJ[4]  (.A(count_8[4]), .B(N_25), .Y(N_26));
    XA1B \count_RNO[3]  (.A(N_24), .B(count_8[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    DFN1 \count[11]  (.D(count_n11), .CLK(GLA), .Q(count_1[11]));
    XA1B \count_RNO[8]  (.A(\count_RNI4LSV[1]_net_1 ), .B(count_1[8]), 
        .C(count_0_sqmuxa_net_1), .Y(N_19));
    NOR2B \count_RNIBDV7[7]  (.A(count_3[7]), .B(count_8[2]), .Y(
        count_n7_0_i_o3_m3_0_a2_0));
    XA1B \count_RNO[5]  (.A(N_26), .B(count_3[5]), .C(
        count_0_sqmuxa_net_1), .Y(N_13));
    XA1B \count_RNO[1]  (.A(count_8[0]), .B(count_8[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    XA1C \count_RNO[11]  (.A(count_1[11]), .B(N_32), .C(
        count_0_sqmuxa_net_1), .Y(count_n11));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_8[2]));
    OR2B \count_RNI3DU7[1]  (.A(count_8[1]), .B(count_8[0]), .Y(N_23));
    GND GND_i (.Y(GND));
    DFN1 \count[9]  (.D(count_n9), .CLK(GLA), .Q(count_1[9]));
    NOR3 \count_RNO[6]  (.A(N_61), .B(count_0_sqmuxa_net_1), .C(N_28), 
        .Y(N_15));
    NOR2 \count_RNO[0]  (.A(count_8[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    OR2A \count_RNO_0[11]  (.A(count_1[10]), .B(N_31), .Y(N_32));
    OR3C count_0_sqmuxa (.A(state1ms_choice_0_dump_start), .B(
        dump_state_0_timer_start), .C(state1ms_choice_0_reset_out), .Y(
        count_0_sqmuxa_net_1));
    NOR2B \count_RNIDLV7[6]  (.A(count_3[5]), .B(count_3[6]), .Y(
        count_n7_0_i_o3_m3_0_a2_2));
    DFN1 \count[6]  (.D(N_15), .CLK(GLA), .Q(count_3[6]));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_8[3]));
    NOR3C \count_RNICKSR[6]  (.A(N_26), .B(count_3[5]), .C(count_3[6]), 
        .Y(N_28));
    OR2B \count_RNITPS31[8]  (.A(count_1[8]), .B(
        \count_RNI4LSV[1]_net_1 ), .Y(N_30));
    NOR2A \count_RNI4LSV[1]  (.A(count_n7_0_i_o3_m3_0_a2_4), .B(N_23), 
        .Y(\count_RNI4LSV[1]_net_1 ));
    OR2 \count_RNO_0[7]  (.A(count_0_sqmuxa_net_1), .B(
        \count_RNI4LSV[1]_net_1 ), .Y(count_n7_0_i_0));
    NOR2B \count_RNI95V7[3]  (.A(count_8[3]), .B(count_8[4]), .Y(
        count_n7_0_i_o3_m3_0_a2_1));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_8[4]));
    DFN1 \count[7]  (.D(N_17), .CLK(GLA), .Q(count_3[7]));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_4(
       count_7,
       GLA,
       state1ms_choice_0_reset_out,
       off_on_state_1_state_over,
       dump_state_0_on_start
    );
output [4:0] count_7;
input  GLA;
input  state1ms_choice_0_reset_out;
input  off_on_state_1_state_over;
input  dump_state_0_on_start;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_14, GND, VCC, GND_0, VCC_0;
    
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_7[0]), .B(count_7[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_7[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_7[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count_7[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    NOR2B \count_RNI08BL[2]  (.A(count_7[2]), .B(N_12), .Y(N_13));
    GND GND_i (.Y(GND));
    NOR2B \count_RNO_0[4]  (.A(count_7[3]), .B(N_13), .Y(N_14));
    XA1B \count_RNO[2]  (.A(N_12), .B(count_7[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(dump_state_0_on_start), .B(
        off_on_state_1_state_over), .C(state1ms_choice_0_reset_out), 
        .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    XA1B \count_RNO[4]  (.A(N_14), .B(count_7[4]), .C(
        count_0_sqmuxa_net_1), .Y(N_11));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_7[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_7[4]));
    NOR2 \count_RNO[0]  (.A(count_7[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    NOR2B \count_RNIVB7E[1]  (.A(count_7[1]), .B(count_7[0]), .Y(N_12));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_7[2]));
    
endmodule


module off_on_coder_4(
       i_6,
       i_7,
       count_7,
       GLA,
       dump_state_0_on_start,
       state1ms_choice_0_reset_out
    );
output [1:1] i_6;
output [0:0] i_7;
input  [4:0] count_7;
input  GLA;
input  dump_state_0_on_start;
input  state1ms_choice_0_reset_out;

    wire \i_0_1[1] , \i_RNO_4[1] , N_17, \i_RNO_5[0] , GND, VCC, GND_0, 
        VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \i_RNO_1[1]  (.A(count_7[1]), .B(count_7[0]), .Y(N_17));
    DFN1 \i[1]  (.D(\i_RNO_4[1] ), .CLK(GLA), .Q(i_6[1]));
    GND GND_i_0 (.Y(GND_0));
    NOR3C \i_RNO[1]  (.A(\i_0_1[1] ), .B(N_17), .C(
        state1ms_choice_0_reset_out), .Y(\i_RNO_4[1] ));
    VCC VCC_i (.Y(VCC));
    NOR3B \i_RNO_0[1]  (.A(count_7[2]), .B(count_7[4]), .C(count_7[3]), 
        .Y(\i_0_1[1] ));
    NOR2B \i_RNO[0]  (.A(state1ms_choice_0_reset_out), .B(
        dump_state_0_on_start), .Y(\i_RNO_5[0] ));
    DFN1 \i[0]  (.D(\i_RNO_5[0] ), .CLK(GLA), .Q(i_7[0]));
    GND GND_i (.Y(GND));
    
endmodule


module DUMP(
       dumpdata,
       dump_cho,
       state1ms_choice_0_dump_start,
       top_code_0_dumpload,
       state1ms_choice_0_bri_cycle,
       bri_div_start_0,
       DUMP_0_dump_off,
       DUMP_0_dump_on,
       state1ms_choice_0_reset_out,
       GLA
    );
input  [11:0] dumpdata;
input  [2:0] dump_cho;
input  state1ms_choice_0_dump_start;
input  top_code_0_dumpload;
input  state1ms_choice_0_bri_cycle;
input  bri_div_start_0;
output DUMP_0_dump_off;
output DUMP_0_dump_on;
input  state1ms_choice_0_reset_out;
input  GLA;

    wire \count_9[0] , \count_9[1] , \count_9[2] , \count_9[3] , 
        \count_9[4] , dump_state_0_off_start, 
        off_on_state_0_state_over, \i_9[0] , \i_8[1] , \i_5[2] , 
        \i_5[3] , \i_1[4] , \i_1[5] , \i_0[6] , \i_0[7] , \i_0[8] , 
        dump_state_0_timer_start, dump_state_0_on_start, \i_7[1] , 
        \i_8[0] , \i_6[1] , \i_7[0] , off_on_state_1_state_over, 
        \count_3[5] , \count_3[6] , \count_3[7] , \count_8[0] , 
        \count_8[1] , \count_8[2] , \count_8[3] , \count_8[4] , 
        \count_1[8] , \count_1[9] , \count_1[10] , \count_1[11] , 
        \count_7[0] , \count_7[1] , \count_7[2] , \count_7[3] , 
        \count_7[4] , GND, VCC, GND_0, VCC_0;
    
    off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_3 
        off_on_timer_0 (.count_9({\count_9[4] , \count_9[3] , 
        \count_9[2] , \count_9[1] , \count_9[0] }), .GLA(GLA), 
        .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out), 
        .dump_state_0_off_start(dump_state_0_off_start), 
        .off_on_state_0_state_over(off_on_state_0_state_over));
    dump_state dump_state_0 (.i_9({\i_9[0] }), .i_8({\i_8[1] }), .i_5({
        \i_5[3] , \i_5[2] }), .i_1({\i_1[5] , \i_1[4] }), .i_0({
        \i_0[8] , \i_0[7] , \i_0[6] }), .dump_state_0_off_start(
        dump_state_0_off_start), .GLA(GLA), 
        .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out), 
        .dump_state_0_timer_start(dump_state_0_timer_start), 
        .dump_state_0_on_start(dump_state_0_on_start));
    off_on_coder_3 off_on_coder_1 (.i_7({\i_7[1] }), .i_8({\i_8[0] }), 
        .count_9({\count_9[4] , \count_9[3] , \count_9[2] , 
        \count_9[1] , \count_9[0] }), .GLA(GLA), 
        .dump_state_0_off_start(dump_state_0_off_start), 
        .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out));
    off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_3 
        off_on_state_1 (.i_6({\i_6[1] }), .i_7({\i_7[0] }), .GLA(GLA), 
        .DUMP_0_dump_on(DUMP_0_dump_on), .off_on_state_1_state_over(
        off_on_state_1_state_over), .state1ms_choice_0_reset_out(
        state1ms_choice_0_reset_out));
    VCC VCC_i_0 (.Y(VCC_0));
    off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_4 
        off_on_state_0 (.i_7({\i_7[1] }), .i_8({\i_8[0] }), .GLA(GLA), 
        .DUMP_0_dump_off(DUMP_0_dump_off), .off_on_state_0_state_over(
        off_on_state_0_state_over), .state1ms_choice_0_reset_out(
        state1ms_choice_0_reset_out));
    dump_coder dump_coder_0 (.i_0({\i_0[8] , \i_0[7] , \i_0[6] }), 
        .i_1({\i_1[5] , \i_1[4] }), .i_5({\i_5[3] , \i_5[2] }), .i_8({
        \i_8[1] }), .i_9({\i_9[0] }), .count_3({\count_3[7] , 
        \count_3[6] , \count_3[5] }), .dump_cho({dump_cho[2], 
        dump_cho[1], dump_cho[0]}), .dumpdata({dumpdata[11], 
        dumpdata[10], dumpdata[9], dumpdata[8], dumpdata[7], 
        dumpdata[6], dumpdata[5], dumpdata[4], dumpdata[3], 
        dumpdata[2], dumpdata[1], dumpdata[0]}), .count_8({
        \count_8[4] , \count_8[3] , \count_8[2] , \count_8[1] , 
        \count_8[0] }), .count_1({\count_1[11] , \count_1[10] , 
        \count_1[9] , \count_1[8] }), .GLA(GLA), .bri_div_start_0(
        bri_div_start_0), .state1ms_choice_0_bri_cycle(
        state1ms_choice_0_bri_cycle), .top_code_0_dumpload(
        top_code_0_dumpload), .state1ms_choice_0_dump_start(
        state1ms_choice_0_dump_start), .state1ms_choice_0_reset_out(
        state1ms_choice_0_reset_out));
    VCC VCC_i (.Y(VCC));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    dump_timer dump_timer_0 (.count_1({\count_1[11] , \count_1[10] , 
        \count_1[9] , \count_1[8] }), .count_8({\count_8[4] , 
        \count_8[3] , \count_8[2] , \count_8[1] , \count_8[0] }), 
        .count_3({\count_3[7] , \count_3[6] , \count_3[5] }), .GLA(GLA)
        , .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out), 
        .dump_state_0_timer_start(dump_state_0_timer_start), 
        .state1ms_choice_0_dump_start(state1ms_choice_0_dump_start));
    off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_4 
        off_on_timer_1 (.count_7({\count_7[4] , \count_7[3] , 
        \count_7[2] , \count_7[1] , \count_7[0] }), .GLA(GLA), 
        .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out), 
        .off_on_state_1_state_over(off_on_state_1_state_over), 
        .dump_state_0_on_start(dump_state_0_on_start));
    off_on_coder_4 off_on_coder_0 (.i_6({\i_6[1] }), .i_7({\i_7[0] }), 
        .count_7({\count_7[4] , \count_7[3] , \count_7[2] , 
        \count_7[1] , \count_7[0] }), .GLA(GLA), 
        .dump_state_0_on_start(dump_state_0_on_start), 
        .state1ms_choice_0_reset_out(state1ms_choice_0_reset_out));
    
endmodule


module long_timer(
       sigtimedata,
       GLA,
       top_code_0_sigrst,
       sigtimeup_c,
       clk_5K,
       net_27
    );
input  [15:0] sigtimedata;
input  GLA;
input  top_code_0_sigrst;
output sigtimeup_c;
input  clk_5K;
input  net_27;

    wire count_n7_0_i_0, \count_RNIS1KE1[1]_net_1 , en_net_1, 
        timeup_0_sqmuxa_13, timeup_0_sqmuxa_2, timeup_0_sqmuxa_1, 
        timeup_0_sqmuxa_10, timeup_0_sqmuxa_12, timeup_0_sqmuxa_0, 
        N_96_i_i_0, timeup_0_sqmuxa_7, timeup_0_sqmuxa_11, N_89_i_i_0, 
        N_101_i_i_0, timeup_0_sqmuxa_6, N_98_i_i_0, N_97_i_i_0, 
        timeup_0_sqmuxa_4, \count[5]_net_1 , N_93_i_i_0, 
        \count[3]_net_1 , N_91_i_i_0, \count[12]_net_1 , N_100_i_i_0, 
        \count[7]_net_1 , N_95_i_i_0, \count[15]_net_1 , N_87_i_i_0, 
        \count[1]_net_1 , clk_5K_en_1_i, count_n7_0_i_o2_m3_0_a2_4, 
        count_n7_0_i_o2_m3_0_a2_1, count_n7_0_i_o2_m3_0_a2_0, 
        count_n7_0_i_o2_m3_0_a2_2, \count[6]_net_1 , \count[4]_net_1 , 
        \count[2]_net_1 , count_n11_0_0_o2_m6_0_a2_7, 
        count_n11_0_0_o2_m6_0_a2_1, N_44_i_0, 
        count_n11_0_0_o2_m6_0_a2_6, count_n11_0_0_o2_m6_0_a2_0, 
        \count[9]_net_1 , \count[10]_net_1 , \count[8]_net_1 , N_5, 
        \count[0]_net_1 , N_7, N_9, N_74, N_11, N_95, N_13, N_96, N_15, 
        N_97, timeup_0_sqmuxa, N_19_i_0, N_17, N_98, 
        \count_RNIAOOQ1[9]_net_1 , count_n10, N_101, count_n11, 
        \count[11]_net_1 , count_n12, N_103, count_n13, N_104, 
        \count[13]_net_1 , count_n9, N_100, count_n0, count_n14, 
        \count[14]_net_1 , N_105, count_n15, N_106, 
        clk_5K_reg1_RNO_net_1, clk_5K_reg1_net_1, clk_5K_reg2_net_1, 
        clk_5K_reg2_RNO_net_1, timeup_RNO_net_1, counte, GND, VCC, 
        GND_0, VCC_0;
    
    XA1A timeup_RNO_9 (.A(\count[3]_net_1 ), .B(sigtimedata[3]), .C(
        N_91_i_i_0), .Y(timeup_0_sqmuxa_6));
    DFN1E1 \count[5]  (.D(N_13), .CLK(GLA), .E(counte), .Q(
        \count[5]_net_1 ));
    XNOR2 timeup_RNO_7 (.A(sigtimedata[2]), .B(\count[2]_net_1 ), .Y(
        N_89_i_i_0));
    DFN1E1 \count[1]  (.D(N_5), .CLK(GLA), .E(counte), .Q(
        \count[1]_net_1 ));
    NOR2B clk_5K_reg1_RNO (.A(net_27), .B(clk_5K), .Y(
        clk_5K_reg1_RNO_net_1));
    NOR3C timeup_RNO_3 (.A(timeup_0_sqmuxa_2), .B(timeup_0_sqmuxa_1), 
        .C(timeup_0_sqmuxa_10), .Y(timeup_0_sqmuxa_13));
    DFN1E1 \count[10]  (.D(count_n10), .CLK(GLA), .E(counte), .Q(
        \count[10]_net_1 ));
    DFN1E1 \count[0]  (.D(count_n0), .CLK(GLA), .E(counte), .Q(
        \count[0]_net_1 ));
    DFN1 clk_5K_reg1 (.D(clk_5K_reg1_RNO_net_1), .CLK(GLA), .Q(
        clk_5K_reg1_net_1));
    DFN1E1 \count[14]  (.D(count_n14), .CLK(GLA), .E(counte), .Q(
        \count[14]_net_1 ));
    NOR3C timeup_RNO_1 (.A(timeup_0_sqmuxa_0), .B(N_96_i_i_0), .C(
        timeup_0_sqmuxa_7), .Y(timeup_0_sqmuxa_12));
    DFN1 timeup (.D(timeup_RNO_net_1), .CLK(GLA), .Q(sigtimeup_c));
    OA1B \count_RNO[7]  (.A(N_98), .B(\count[7]_net_1 ), .C(
        count_n7_0_i_0), .Y(N_17));
    XA1C \count_RNO[15]  (.A(\count[15]_net_1 ), .B(N_106), .C(
        en_net_1), .Y(count_n15));
    NOR2B \count_RNIN0LB[7]  (.A(\count[7]_net_1 ), .B(
        \count[8]_net_1 ), .Y(count_n11_0_0_o2_m6_0_a2_0));
    NOR2A clk_5K_reg2_RNILRUA (.A(clk_5K_reg1_net_1), .B(
        clk_5K_reg2_net_1), .Y(clk_5K_en_1_i));
    NOR2B \count_RNI71V21[5]  (.A(\count[5]_net_1 ), .B(N_96), .Y(N_97)
        );
    XA1A timeup_RNO_6 (.A(\count[5]_net_1 ), .B(sigtimedata[5]), .C(
        N_93_i_i_0), .Y(timeup_0_sqmuxa_7));
    XA1B \count_RNO[2]  (.A(N_44_i_0), .B(\count[2]_net_1 ), .C(
        en_net_1), .Y(N_7));
    XA1C \count_RNO[9]  (.A(N_100), .B(\count[9]_net_1 ), .C(en_net_1), 
        .Y(count_n9));
    AO1A timeup_RNIANVP (.A(sigtimeup_c), .B(clk_5K_en_1_i), .C(
        en_net_1), .Y(counte));
    OR2A \count_RNO_0[10]  (.A(\count[9]_net_1 ), .B(N_100), .Y(N_101));
    VCC VCC_i (.Y(VCC));
    XA1B \count_RNO[4]  (.A(N_95), .B(\count[4]_net_1 ), .C(en_net_1), 
        .Y(N_11));
    DFN1E1 \count[8]  (.D(N_19_i_0), .CLK(GLA), .E(counte), .Q(
        \count[8]_net_1 ));
    XA1A timeup_RNO_19 (.A(\count[12]_net_1 ), .B(sigtimedata[12]), .C(
        N_100_i_i_0), .Y(timeup_0_sqmuxa_4));
    NOR3C timeup_RNO_12 (.A(N_98_i_i_0), .B(N_97_i_i_0), .C(
        timeup_0_sqmuxa_4), .Y(timeup_0_sqmuxa_10));
    XNOR2 timeup_RNO_16 (.A(sigtimedata[0]), .B(\count[0]_net_1 ), .Y(
        N_87_i_i_0));
    XA1A timeup_RNO_10 (.A(\count[7]_net_1 ), .B(sigtimedata[7]), .C(
        N_95_i_i_0), .Y(timeup_0_sqmuxa_2));
    XA1C \count_RNO[10]  (.A(N_101), .B(\count[10]_net_1 ), .C(
        en_net_1), .Y(count_n10));
    NOR2B \count_RNI90LB[1]  (.A(\count[1]_net_1 ), .B(
        \count[0]_net_1 ), .Y(N_44_i_0));
    DFN1E1 \count[15]  (.D(count_n15), .CLK(GLA), .E(counte), .Q(
        \count[15]_net_1 ));
    XA1B \count_RNO[3]  (.A(N_74), .B(\count[3]_net_1 ), .C(en_net_1), 
        .Y(N_9));
    OR2A \count_RNINFOR1[12]  (.A(\count[12]_net_1 ), .B(N_103), .Y(
        N_104));
    DFN1E1 \count[11]  (.D(count_n11), .CLK(GLA), .E(counte), .Q(
        \count[11]_net_1 ));
    XNOR2 timeup_RNO_15 (.A(sigtimedata[8]), .B(\count[8]_net_1 ), .Y(
        N_95_i_i_0));
    XA1C \count_RNO[8]  (.A(\count[8]_net_1 ), .B(
        \count_RNIS1KE1[1]_net_1 ), .C(en_net_1), .Y(N_19_i_0));
    NOR2B \count_RNIR5A6[10]  (.A(\count[10]_net_1 ), .B(
        \count[2]_net_1 ), .Y(count_n11_0_0_o2_m6_0_a2_1));
    XNOR2 timeup_RNO_18 (.A(sigtimedata[10]), .B(\count[10]_net_1 ), 
        .Y(N_97_i_i_0));
    NOR2B \count_RNIF0LB[3]  (.A(\count[3]_net_1 ), .B(
        \count[4]_net_1 ), .Y(count_n7_0_i_o2_m3_0_a2_1));
    NOR2B \count_RNIUG4T[4]  (.A(\count[4]_net_1 ), .B(N_95), .Y(N_96));
    DFN1E1 \count[13]  (.D(count_n13), .CLK(GLA), .E(counte), .Q(
        \count[13]_net_1 ));
    XA1B \count_RNO[5]  (.A(N_96), .B(\count[5]_net_1 ), .C(en_net_1), 
        .Y(N_13));
    XA1B \count_RNO[1]  (.A(\count[0]_net_1 ), .B(\count[1]_net_1 ), 
        .C(en_net_1), .Y(N_5));
    XA1C \count_RNO[11]  (.A(\count[11]_net_1 ), .B(
        \count_RNIAOOQ1[9]_net_1 ), .C(en_net_1), .Y(count_n11));
    OR2A \count_RNO_1[7]  (.A(\count_RNIS1KE1[1]_net_1 ), .B(en_net_1), 
        .Y(count_n7_0_i_0));
    OR2A \count_RNIFH8S1[13]  (.A(\count[13]_net_1 ), .B(N_104), .Y(
        N_105));
    NOR2B clk_5K_reg2_RNO (.A(net_27), .B(clk_5K_reg1_net_1), .Y(
        clk_5K_reg2_RNO_net_1));
    DFN1E1 \count[2]  (.D(N_7), .CLK(GLA), .E(counte), .Q(
        \count[2]_net_1 ));
    OR2B en (.A(top_code_0_sigrst), .B(net_27), .Y(en_net_1));
    OR2B \count_RNIAOOQ1[9]  (.A(count_n11_0_0_o2_m6_0_a2_7), .B(
        count_n11_0_0_o2_m6_0_a2_6), .Y(\count_RNIAOOQ1[9]_net_1 ));
    NOR2B \count_RNIFGFH[2]  (.A(\count[2]_net_1 ), .B(N_44_i_0), .Y(
        N_74));
    GND GND_i (.Y(GND));
    OR2B \count_RNIS1KE1[1]  (.A(count_n7_0_i_o2_m3_0_a2_4), .B(
        N_44_i_0), .Y(\count_RNIS1KE1[1]_net_1 ));
    DFN1E1 \count[9]  (.D(count_n9), .CLK(GLA), .E(counte), .Q(
        \count[9]_net_1 ));
    XA1B \count_RNO[6]  (.A(N_97), .B(\count[6]_net_1 ), .C(en_net_1), 
        .Y(N_15));
    XA1C \count_RNO[12]  (.A(N_103), .B(\count[12]_net_1 ), .C(
        en_net_1), .Y(count_n12));
    NOR2 \count_RNO[0]  (.A(en_net_1), .B(\count[0]_net_1 ), .Y(
        count_n0));
    XNOR2 timeup_RNO_14 (.A(sigtimedata[4]), .B(\count[4]_net_1 ), .Y(
        N_91_i_i_0));
    NOR3C \count_RNIJ6KT[10]  (.A(count_n7_0_i_o2_m3_0_a2_1), .B(
        count_n11_0_0_o2_m6_0_a2_1), .C(N_44_i_0), .Y(
        count_n11_0_0_o2_m6_0_a2_7));
    XNOR2 timeup_RNO_17 (.A(sigtimedata[11]), .B(\count[11]_net_1 ), 
        .Y(N_98_i_i_0));
    NOR3C timeup_RNO_0 (.A(timeup_0_sqmuxa_12), .B(timeup_0_sqmuxa_11), 
        .C(timeup_0_sqmuxa_13), .Y(timeup_0_sqmuxa));
    DFN1E1 \count[6]  (.D(N_15), .CLK(GLA), .E(counte), .Q(
        \count[6]_net_1 ));
    NOR3C timeup_RNO_2 (.A(N_89_i_i_0), .B(N_101_i_i_0), .C(
        timeup_0_sqmuxa_6), .Y(timeup_0_sqmuxa_11));
    XNOR2 timeup_RNO_13 (.A(sigtimedata[6]), .B(\count[6]_net_1 ), .Y(
        N_93_i_i_0));
    DFN1E1 \count[3]  (.D(N_9), .CLK(GLA), .E(counte), .Q(
        \count[3]_net_1 ));
    OR2A \count_RNI8IEK1[8]  (.A(\count[8]_net_1 ), .B(
        \count_RNIS1KE1[1]_net_1 ), .Y(N_100));
    XA1A timeup_RNO_11 (.A(\count[15]_net_1 ), .B(sigtimedata[15]), .C(
        N_87_i_i_0), .Y(timeup_0_sqmuxa_1));
    NOR3C \count_RNIJ1V21[7]  (.A(count_n7_0_i_o2_m3_0_a2_1), .B(
        count_n7_0_i_o2_m3_0_a2_0), .C(count_n7_0_i_o2_m3_0_a2_2), .Y(
        count_n7_0_i_o2_m3_0_a2_4));
    XA1C \count_RNO[14]  (.A(\count[14]_net_1 ), .B(N_105), .C(
        en_net_1), .Y(count_n14));
    NOR2B \count_RNIH0LB[7]  (.A(\count[7]_net_1 ), .B(
        \count[2]_net_1 ), .Y(count_n7_0_i_o2_m3_0_a2_0));
    XA1C \count_RNO[13]  (.A(N_104), .B(\count[13]_net_1 ), .C(
        en_net_1), .Y(count_n13));
    NOR2B \count_RNO_0[7]  (.A(\count[6]_net_1 ), .B(N_97), .Y(N_98));
    DFN1 clk_5K_reg2 (.D(clk_5K_reg2_RNO_net_1), .CLK(GLA), .Q(
        clk_5K_reg2_net_1));
    XNOR2 timeup_RNO_8 (.A(sigtimedata[14]), .B(\count[14]_net_1 ), .Y(
        N_101_i_i_0));
    NOR2B \count_RNIJ0LB[5]  (.A(\count[5]_net_1 ), .B(
        \count[6]_net_1 ), .Y(count_n7_0_i_o2_m3_0_a2_2));
    XNOR2 timeup_RNO_20 (.A(sigtimedata[13]), .B(\count[13]_net_1 ), 
        .Y(N_100_i_i_0));
    OR2A \count_RNO_0[15]  (.A(\count[14]_net_1 ), .B(N_105), .Y(N_106)
        );
    NOR2B \count_RNIM0AN[3]  (.A(\count[3]_net_1 ), .B(N_74), .Y(N_95));
    OA1B timeup_RNO (.A(timeup_0_sqmuxa), .B(sigtimeup_c), .C(en_net_1)
        , .Y(timeup_RNO_net_1));
    DFN1E1 \count[4]  (.D(N_11), .CLK(GLA), .E(counte), .Q(
        \count[4]_net_1 ));
    OR2A \count_RNI0I8R1[11]  (.A(\count[11]_net_1 ), .B(
        \count_RNIAOOQ1[9]_net_1 ), .Y(N_103));
    XA1A timeup_RNO_4 (.A(\count[1]_net_1 ), .B(sigtimedata[1]), .C(
        clk_5K_en_1_i), .Y(timeup_0_sqmuxa_0));
    DFN1E1 \count[12]  (.D(count_n12), .CLK(GLA), .E(counte), .Q(
        \count[12]_net_1 ));
    NOR3C \count_RNINH4T[9]  (.A(count_n11_0_0_o2_m6_0_a2_0), .B(
        \count[9]_net_1 ), .C(count_n7_0_i_o2_m3_0_a2_2), .Y(
        count_n11_0_0_o2_m6_0_a2_6));
    DFN1E1 \count[7]  (.D(N_17), .CLK(GLA), .E(counte), .Q(
        \count[7]_net_1 ));
    XNOR2 timeup_RNO_5 (.A(sigtimedata[9]), .B(\count[9]_net_1 ), .Y(
        N_96_i_i_0));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module clk_div500(
       GLA,
       pllclk_0_GLB,
       net_27,
       clk_5K
    );
input  GLA;
input  pllclk_0_GLB;
input  net_27;
output clk_5K;

    wire \DWACT_ADD_CI_0_g_array_2[0] , \DWACT_ADD_CI_0_g_array_1[0] , 
        \DWACT_ADD_CI_0_pog_array_1[0] , \DWACT_ADD_CI_0_g_array_3[0] , 
        \DWACT_ADD_CI_0_pog_array_2[0] , \DWACT_ADD_CI_0_TMP[0] , 
        \count[1]_net_1 , \DWACT_ADD_CI_0_g_array_11[0] , 
        \DWACT_ADD_CI_0_pog_array_1_1[0] , 
        \DWACT_ADD_CI_0_g_array_12_1[0] , \count[4]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12[0] , \count[2]_net_1 , 
        \DWACT_ADD_CI_0_g_array_12_2[0] , \count[6]_net_1 , 
        count_0_sqmuxa_6, clk_5M_en, \count[0]_net_1 , 
        count_0_sqmuxa_5, \count[5]_net_1 , count_0_sqmuxa_2, 
        count_0_sqmuxa_4, \count[8]_net_1 , \count[3]_net_1 , 
        \count[7]_net_1 , count_0_sqmuxa, N_41, clk_5M_reg1_net_1, 
        clk_5M_reg2_net_1, \count_5[1] , I_32, \count_5[2] , I_35, 
        \count_5[3] , I_37, \count_5[4] , I_30, \count_5[5] , I_33, 
        \count_5[6] , I_36, \count_5[7] , I_38_0, \count_5[8] , I_34, 
        \count_5[0] , \DWACT_ADD_CI_0_partial_sum[0] , 
        clk_5K_RNO_net_1, clk_5M_reg2_RNO_net_1, clk_5M_reg1_RNO_net_1, 
        \DWACT_ADD_CI_0_pog_array_1_2[0] , GND, VCC, GND_0, VCC_0;
    
    XOR2 un1_count_1_I_37 (.A(\count[3]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12[0] ), .Y(I_37));
    DFN1 \count[5]  (.D(\count_5[5] ), .CLK(GLA), .Q(\count[5]_net_1 ));
    NOR2A clk_5M_reg2_RNI74E6 (.A(clk_5M_reg1_net_1), .B(
        clk_5M_reg2_net_1), .Y(clk_5M_en));
    NOR2B un1_count_1_I_47 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \count[4]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_1[0] ));
    NOR2B clk_5M_reg2_RNO (.A(net_27), .B(clk_5M_reg1_net_1), .Y(
        clk_5M_reg2_RNO_net_1));
    DFN1 \count[1]  (.D(\count_5[1] ), .CLK(GLA), .Q(\count[1]_net_1 ));
    NOR2B un1_count_1_I_49 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \count[2]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12[0] ));
    DFN1 \count[0]  (.D(\count_5[0] ), .CLK(GLA), .Q(\count[0]_net_1 ));
    AND2 un1_count_1_I_1 (.A(\count[0]_net_1 ), .B(clk_5M_en), .Y(
        \DWACT_ADD_CI_0_TMP[0] ));
    AND2 un1_count_1_I_52 (.A(\count[2]_net_1 ), .B(\count[3]_net_1 ), 
        .Y(\DWACT_ADD_CI_0_pog_array_1[0] ));
    NOR3B \count_RNO[7]  (.A(net_27), .B(I_38_0), .C(count_0_sqmuxa), 
        .Y(\count_5[7] ));
    DFN1 clk_5M_reg2 (.D(clk_5M_reg2_RNO_net_1), .CLK(GLA), .Q(
        clk_5M_reg2_net_1));
    NOR3B \count_RNO[2]  (.A(net_27), .B(I_35), .C(count_0_sqmuxa), .Y(
        \count_5[2] ));
    AND2 un1_count_1_I_53 (.A(\count[4]_net_1 ), .B(\count[5]_net_1 ), 
        .Y(\DWACT_ADD_CI_0_pog_array_1_1[0] ));
    VCC VCC_i (.Y(VCC));
    NOR3B \count_RNO[4]  (.A(net_27), .B(I_30), .C(count_0_sqmuxa), .Y(
        \count_5[4] ));
    DFN1 \count[8]  (.D(\count_5[8] ), .CLK(GLA), .Q(\count[8]_net_1 ));
    NOR2B un1_count_1_I_50 (.A(\DWACT_ADD_CI_0_g_array_11[0] ), .B(
        \count[6]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_12_2[0] ));
    NOR3B \count_RNO[3]  (.A(net_27), .B(I_37), .C(count_0_sqmuxa), .Y(
        \count_5[3] ));
    NOR3B \count_RNO[8]  (.A(net_27), .B(I_34), .C(count_0_sqmuxa), .Y(
        \count_5[8] ));
    AND2 un1_count_1_I_54 (.A(\count[6]_net_1 ), .B(\count[7]_net_1 ), 
        .Y(\DWACT_ADD_CI_0_pog_array_1_2[0] ));
    DFN1 clk_5M_reg1 (.D(clk_5M_reg1_RNO_net_1), .CLK(GLA), .Q(
        clk_5M_reg1_net_1));
    NOR3B \count_RNO[5]  (.A(net_27), .B(I_33), .C(count_0_sqmuxa), .Y(
        \count_5[5] ));
    NOR3B \count_RNO[1]  (.A(net_27), .B(I_32), .C(count_0_sqmuxa), .Y(
        \count_5[1] ));
    XOR2 un1_count_1_I_36 (.A(\count[6]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_11[0] ), .Y(I_36));
    DFN1 \count[2]  (.D(\count_5[2] ), .CLK(GLA), .Q(\count[2]_net_1 ));
    NOR2B un1_count_1_I_46 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_2[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_3[0] ));
    XOR2 un1_count_1_I_32 (.A(\count[1]_net_1 ), .B(
        \DWACT_ADD_CI_0_TMP[0] ), .Y(I_32));
    NOR3A \count_RNIA69L[0]  (.A(clk_5M_en), .B(\count[1]_net_1 ), .C(
        \count[0]_net_1 ), .Y(count_0_sqmuxa_6));
    GND GND_i (.Y(GND));
    NOR3B \count_RNO[6]  (.A(net_27), .B(I_36), .C(count_0_sqmuxa), .Y(
        \count_5[6] ));
    OR3A \count_RNO[0]  (.A(net_27), .B(count_0_sqmuxa), .C(
        \DWACT_ADD_CI_0_partial_sum[0] ), .Y(\count_5[0] ));
    XOR2 un1_count_1_I_33 (.A(\count[5]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_1[0] ), .Y(I_33));
    NOR2B un1_count_1_I_43 (.A(\DWACT_ADD_CI_0_g_array_2[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_11[0] ));
    NOR2B \count_RNIF2RE[7]  (.A(\count[6]_net_1 ), .B(
        \count[7]_net_1 ), .Y(count_0_sqmuxa_2));
    NOR2B clk_5M_reg1_RNO (.A(net_27), .B(pllclk_0_GLB), .Y(
        clk_5M_reg1_RNO_net_1));
    XOR2 un1_count_1_I_30 (.A(\count[4]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_2[0] ), .Y(I_30));
    NOR2B un1_count_1_I_40 (.A(\DWACT_ADD_CI_0_TMP[0] ), .B(
        \count[1]_net_1 ), .Y(\DWACT_ADD_CI_0_g_array_1[0] ));
    DFN1 \count[6]  (.D(\count_5[6] ), .CLK(GLA), .Q(\count[6]_net_1 ));
    XOR2 un1_count_1_I_21 (.A(\count[0]_net_1 ), .B(clk_5M_en), .Y(
        \DWACT_ADD_CI_0_partial_sum[0] ));
    DFN1 \count[3]  (.D(\count_5[3] ), .CLK(GLA), .Q(\count[3]_net_1 ));
    MX2B clk_5K_RNO_0 (.A(clk_5K), .B(clk_5K), .S(count_0_sqmuxa), .Y(
        N_41));
    NOR2B clk_5K_RNO (.A(net_27), .B(N_41), .Y(clk_5K_RNO_net_1));
    AND2 un1_count_1_I_51 (.A(\DWACT_ADD_CI_0_pog_array_1_1[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1_2[0] ), .Y(
        \DWACT_ADD_CI_0_pog_array_2[0] ));
    XOR2 un1_count_1_I_34 (.A(\count[8]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_3[0] ), .Y(I_34));
    NOR2B un1_count_1_I_44 (.A(\DWACT_ADD_CI_0_g_array_1[0] ), .B(
        \DWACT_ADD_CI_0_pog_array_1[0] ), .Y(
        \DWACT_ADD_CI_0_g_array_2[0] ));
    XOR2 un1_count_1_I_35 (.A(\count[2]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_1[0] ), .Y(I_35));
    XOR2 un1_count_1_I_38 (.A(\count[7]_net_1 ), .B(
        \DWACT_ADD_CI_0_g_array_12_2[0] ), .Y(I_38_0));
    NOR3C \count_RNIQ4MT[5]  (.A(\count[5]_net_1 ), .B(
        \count[4]_net_1 ), .C(count_0_sqmuxa_2), .Y(count_0_sqmuxa_5));
    DFN1 clk_5K_inst_1 (.D(clk_5K_RNO_net_1), .CLK(GLA), .Q(clk_5K));
    DFN1 \count[4]  (.D(\count_5[4] ), .CLK(GLA), .Q(\count[4]_net_1 ));
    DFN1 \count[7]  (.D(\count_5[7] ), .CLK(GLA), .Q(\count[7]_net_1 ));
    NOR3C \count_RNIKU792[0]  (.A(count_0_sqmuxa_5), .B(
        count_0_sqmuxa_4), .C(count_0_sqmuxa_6), .Y(count_0_sqmuxa));
    NOR3B \count_RNIGJ8M[8]  (.A(\count[2]_net_1 ), .B(
        \count[8]_net_1 ), .C(\count[3]_net_1 ), .Y(count_0_sqmuxa_4));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module pllclk(
       pllclk_VCC,
       pllclk_GND,
       OCX40MHz_c,
       pllclk_0_GLB,
       GLA
    );
input  pllclk_VCC;
input  pllclk_GND;
input  OCX40MHz_c;
output pllclk_0_GLB;
output GLA;

    wire Core_GLC, Core_LOCK, Core_YB, Core_YC, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    PLL #( .VCOFREQUENCY(100.000000) )  Core (.CLKA(OCX40MHz_c), 
        .EXTFB(pllclk_GND), .POWERDOWN(pllclk_VCC), .GLA(GLA), .LOCK(
        Core_LOCK), .GLB(pllclk_0_GLB), .YB(Core_YB), .GLC(Core_GLC), 
        .YC(Core_YC), .OADIV0(pllclk_GND), .OADIV1(pllclk_GND), 
        .OADIV2(pllclk_GND), .OADIV3(pllclk_GND), .OADIV4(pllclk_GND), 
        .OAMUX0(pllclk_GND), .OAMUX1(pllclk_GND), .OAMUX2(pllclk_VCC), 
        .DLYGLA0(pllclk_GND), .DLYGLA1(pllclk_GND), .DLYGLA2(
        pllclk_GND), .DLYGLA3(pllclk_GND), .DLYGLA4(pllclk_GND), 
        .OBDIV0(pllclk_VCC), .OBDIV1(pllclk_VCC), .OBDIV2(pllclk_GND), 
        .OBDIV3(pllclk_GND), .OBDIV4(pllclk_VCC), .OBMUX0(pllclk_GND), 
        .OBMUX1(pllclk_VCC), .OBMUX2(pllclk_GND), .DLYYB0(pllclk_GND), 
        .DLYYB1(pllclk_GND), .DLYYB2(pllclk_GND), .DLYYB3(pllclk_GND), 
        .DLYYB4(pllclk_GND), .DLYGLB0(pllclk_GND), .DLYGLB1(pllclk_GND)
        , .DLYGLB2(pllclk_GND), .DLYGLB3(pllclk_GND), .DLYGLB4(
        pllclk_GND), .OCDIV0(pllclk_GND), .OCDIV1(pllclk_GND), .OCDIV2(
        pllclk_GND), .OCDIV3(pllclk_GND), .OCDIV4(pllclk_GND), .OCMUX0(
        pllclk_GND), .OCMUX1(pllclk_GND), .OCMUX2(pllclk_GND), .DLYYC0(
        pllclk_GND), .DLYYC1(pllclk_GND), .DLYYC2(pllclk_GND), .DLYYC3(
        pllclk_GND), .DLYYC4(pllclk_GND), .DLYGLC0(pllclk_GND), 
        .DLYGLC1(pllclk_GND), .DLYGLC2(pllclk_GND), .DLYGLC3(
        pllclk_GND), .DLYGLC4(pllclk_GND), .FINDIV0(pllclk_VCC), 
        .FINDIV1(pllclk_VCC), .FINDIV2(pllclk_VCC), .FINDIV3(
        pllclk_GND), .FINDIV4(pllclk_GND), .FINDIV5(pllclk_GND), 
        .FINDIV6(pllclk_GND), .FBDIV0(pllclk_VCC), .FBDIV1(pllclk_VCC), 
        .FBDIV2(pllclk_GND), .FBDIV3(pllclk_GND), .FBDIV4(pllclk_VCC), 
        .FBDIV5(pllclk_GND), .FBDIV6(pllclk_GND), .FBDLY0(pllclk_GND), 
        .FBDLY1(pllclk_GND), .FBDLY2(pllclk_GND), .FBDLY3(pllclk_GND), 
        .FBDLY4(pllclk_GND), .FBSEL0(pllclk_VCC), .FBSEL1(pllclk_GND), 
        .XDLYSEL(pllclk_GND), .VCOSEL0(pllclk_GND), .VCOSEL1(
        pllclk_GND), .VCOSEL2(pllclk_VCC));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module ClockManagement(
       sigtimedata,
       OCX40MHz_c,
       ClockManagement_GND,
       ClockManagement_VCC,
       net_27,
       clk_5K,
       sigtimeup_c,
       top_code_0_sigrst,
       GLA
    );
input  [15:0] sigtimedata;
input  OCX40MHz_c;
input  ClockManagement_GND;
input  ClockManagement_VCC;
input  net_27;
output clk_5K;
output sigtimeup_c;
input  top_code_0_sigrst;
output GLA;

    wire pllclk_0_GLB, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    long_timer long_timer_0 (.sigtimedata({sigtimedata[15], 
        sigtimedata[14], sigtimedata[13], sigtimedata[12], 
        sigtimedata[11], sigtimedata[10], sigtimedata[9], 
        sigtimedata[8], sigtimedata[7], sigtimedata[6], sigtimedata[5], 
        sigtimedata[4], sigtimedata[3], sigtimedata[2], sigtimedata[1], 
        sigtimedata[0]}), .GLA(GLA), .top_code_0_sigrst(
        top_code_0_sigrst), .sigtimeup_c(sigtimeup_c), .clk_5K(clk_5K), 
        .net_27(net_27));
    clk_div500 clk_div500_0 (.GLA(GLA), .pllclk_0_GLB(pllclk_0_GLB), 
        .net_27(net_27), .clk_5K(clk_5K));
    GND GND_i_0 (.Y(GND_0));
    pllclk pllclk_0 (.pllclk_VCC(ClockManagement_VCC), .pllclk_GND(
        ClockManagement_GND), .OCX40MHz_c(OCX40MHz_c), .pllclk_0_GLB(
        pllclk_0_GLB), .GLA(GLA));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module pd_pluse_coder(
       i_0,
       i_4,
       i_5,
       pd_pluse_data,
       i_0_0_0,
       pd_pluse_choice,
       count_0,
       count_2,
       count_5,
       ddsclkout_c,
       GLA,
       bri_dump_sw_0_tetw_pluse,
       net_51,
       pulse_start_c,
       top_code_0_pd_pluse_load,
       net_27
    );
output [5:4] i_0;
output [3:2] i_4;
output [0:0] i_5;
input  [15:0] pd_pluse_data;
output i_0_0_0;
input  [3:0] pd_pluse_choice;
input  [15:8] count_0;
input  [7:5] count_2;
input  [4:0] count_5;
input  ddsclkout_c;
input  GLA;
input  bri_dump_sw_0_tetw_pluse;
input  net_51;
input  pulse_start_c;
input  top_code_0_pd_pluse_load;
input  net_27;

    wire \i_0_15[4] , \i_0_12[4] , \i_0_11[4] , \i_0_13[4] , 
        \i_0_2[4] , \i_0_1[4] , \i_0_10[4] , \un1_count_1_0_0_i_0[0] , 
        \un1_count_1_12_i_0[0] , \i_0_8[4] , \un1_count_1_4_i_0[0] , 
        \un1_count_1_1_i_0[0] , \i_0_6[4] , \un1_count_1_7_i_0[0] , 
        \un1_count_1_5_i_0[0] , \i_0_4[4] , \pd_pluse_data3[3]_net_1 , 
        \i_0_0[4] , \pd_pluse_data3[6]_net_1 , \un1_count_1_9_i_0[0] , 
        \pd_pluse_data3[10]_net_1 , \un1_count_1_13_i_0[0] , 
        \pd_pluse_data3[14]_net_1 , \un1_count_1_2_i_0[0] , 
        \pd_pluse_data3[8]_net_1 , \un1_count_1_11_i_0[0] , 
        \pd_pluse_data3[15]_net_1 , \i_reg10_NE_13[0] , 
        \i_reg10_NE_5[0] , \i_reg10_NE_4[0] , \i_reg10_NE_11[0] , 
        \i_reg10_NE_12[0] , \i_reg10_NE_1[0] , \i_reg10_NE_0[0] , 
        \i_reg10_NE_9[0] , \i_reg10_12_i[0] , \i_reg10_9_i[0] , 
        \i_reg10_NE_7[0] , \i_reg10_5_i[0] , \i_reg10_2_i[0] , 
        \i_reg10_NE_3[0] , \pd_pluse_data1[0]_net_1 , \i_reg10_3_i[0] , 
        \pd_pluse_data1[4]_net_1 , \i_reg10_6_i[0] , 
        \pd_pluse_data1[13]_net_1 , \i_reg10_1_i[0] , 
        \pd_pluse_data1[7]_net_1 , \i_reg10_10_i[0] , 
        \pd_pluse_data1[11]_net_1 , \i_reg10_14_i[0] , 
        \pd_pluse_data1[15]_net_1 , \i_reg10_8_i[0] , 
        \un1_count_NE_12[0] , \un1_count_NE_3[0] , \un1_count_NE_2[0] , 
        \un1_count_NE_8[0] , \un1_count_NE_11[0] , \un1_count_12_i[0] , 
        \un1_count_9_i[0] , \un1_count_NE_7[0] , \un1_count_NE_10[0] , 
        \un1_count_1_0_i[0] , \un1_count_13_i[0] , \un1_count_NE_5[0] , 
        \un1_count_8_i[0] , \un1_count_15_i[0] , \un1_count_NE_1[0] , 
        \pd_pluse_data2[0]_net_1 , \un1_count_3_i[0] , 
        \pd_pluse_data2[4]_net_1 , \un1_count_6_i[0] , 
        \pd_pluse_data2[7]_net_1 , \un1_count_10_i[0] , 
        \pd_pluse_data2[2]_net_1 , \un1_count_5_i[0] , 
        \pd_pluse_data2[11]_net_1 , \un1_count_14_i[0] , N_12, 
        \i_RNO_2[3] , \un1_count_i_i_0[0] , \i_reg10_NE[0] , 
        \i_RNO_0[4]_net_1 , pd_pluse_data1_0_sqmuxa, 
        pd_pluse_data2_1_sqmuxa, pd_pluse_data3_1_sqmuxa, 
        \pd_pluse_data2[15]_net_1 , \pd_pluse_data1[14]_net_1 , 
        \pd_pluse_data2[14]_net_1 , \pd_pluse_data2[13]_net_1 , 
        \pd_pluse_data3[13]_net_1 , \pd_pluse_data1[12]_net_1 , 
        \pd_pluse_data2[12]_net_1 , \pd_pluse_data3[12]_net_1 , 
        \pd_pluse_data3[11]_net_1 , \pd_pluse_data1[10]_net_1 , 
        \pd_pluse_data2[10]_net_1 , \pd_pluse_data1[9]_net_1 , 
        \pd_pluse_data2[9]_net_1 , \pd_pluse_data3[9]_net_1 , 
        \pd_pluse_data1[8]_net_1 , \pd_pluse_data2[8]_net_1 , 
        \pd_pluse_data3[7]_net_1 , \pd_pluse_data1[6]_net_1 , 
        \pd_pluse_data2[6]_net_1 , \pd_pluse_data1[5]_net_1 , 
        \pd_pluse_data2[5]_net_1 , \pd_pluse_data3[5]_net_1 , 
        \pd_pluse_data3[4]_net_1 , \pd_pluse_data1[3]_net_1 , 
        \pd_pluse_data2[3]_net_1 , \pd_pluse_data1[2]_net_1 , 
        \pd_pluse_data3[2]_net_1 , \pd_pluse_data1[1]_net_1 , 
        \pd_pluse_data2[1]_net_1 , \pd_pluse_data3[1]_net_1 , 
        \pd_pluse_data3[0]_net_1 , \i_RNO_2[0] , \i_RNO_2[2] , 
        \i_RNO_0[5] , GND, VCC, GND_0, VCC_0;
    
    XA1A \pd_pluse_data1_RNIO6BI[15]  (.A(\pd_pluse_data1[15]_net_1 ), 
        .B(count_0[15]), .C(\i_reg10_8_i[0] ), .Y(\i_reg10_NE_0[0] ));
    NOR3C \pd_pluse_data1_RNI89791[2]  (.A(\i_reg10_5_i[0] ), .B(
        \i_reg10_2_i[0] ), .C(\i_reg10_NE_3[0] ), .Y(\i_reg10_NE_9[0] )
        );
    NOR3B pd_pluse_data1_0_sqmuxa_0_a2 (.A(pd_pluse_choice[0]), .B(
        N_12), .C(pd_pluse_choice[1]), .Y(pd_pluse_data1_0_sqmuxa));
    DFN1E1 \pd_pluse_data3[9]  (.D(pd_pluse_data[9]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[9]_net_1 ));
    XA1A \pd_pluse_data2_RNIQPND[11]  (.A(\pd_pluse_data2[11]_net_1 ), 
        .B(count_0[11]), .C(\un1_count_14_i[0] ), .Y(
        \un1_count_NE_1[0] ));
    DFN1E1 \pd_pluse_data2[14]  (.D(pd_pluse_data[14]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[14]_net_1 ));
    XNOR2 \pd_pluse_data2_RNIOVEB[8]  (.A(count_0[8]), .B(
        \pd_pluse_data2[8]_net_1 ), .Y(\un1_count_8_i[0] ));
    XA1A \i_RNO_11[4]  (.A(\pd_pluse_data3[8]_net_1 ), .B(count_0[8]), 
        .C(\un1_count_1_11_i_0[0] ), .Y(\i_0_1[4] ));
    DFN1E1 \pd_pluse_data3[0]  (.D(pd_pluse_data[0]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[0]_net_1 ));
    NOR3B \i_RNO[4]  (.A(\i_0_15[4] ), .B(\i_reg10_NE[0] ), .C(
        \un1_count_i_i_0[0] ), .Y(\i_RNO_0[4]_net_1 ));
    DFN1E1 \pd_pluse_data2[15]  (.D(pd_pluse_data[15]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[15]_net_1 ));
    DFN1 \i[2]  (.D(\i_RNO_2[2] ), .CLK(ddsclkout_c), .Q(i_4[2]));
    NOR3C \i_RNO[3]  (.A(\un1_count_i_i_0[0] ), .B(net_27), .C(
        \i_reg10_NE[0] ), .Y(\i_RNO_2[3] ));
    DFN1E1 \pd_pluse_data2[11]  (.D(pd_pluse_data[11]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[11]_net_1 ));
    XNOR2 \pd_pluse_data1_RNIRQR6[12]  (.A(count_0[12]), .B(
        \pd_pluse_data1[12]_net_1 ), .Y(\i_reg10_12_i[0] ));
    XA1A \pd_pluse_data1_RNIOPND[11]  (.A(\pd_pluse_data1[11]_net_1 ), 
        .B(count_0[11]), .C(\i_reg10_14_i[0] ), .Y(\i_reg10_NE_1[0] ));
    DFN1E1 \pd_pluse_data3[6]  (.D(pd_pluse_data[6]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[6]_net_1 ));
    DFN1E1 \pd_pluse_data1[10]  (.D(pd_pluse_data[10]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[10]_net_1 ));
    XNOR2 \pd_pluse_data2_RNISQR6[12]  (.A(count_0[12]), .B(
        \pd_pluse_data2[12]_net_1 ), .Y(\un1_count_12_i[0] ));
    NOR2B \i_0[1]  (.A(net_51), .B(net_27), .Y(i_0_0_0));
    DFN1 \i[3]  (.D(\i_RNO_2[3] ), .CLK(ddsclkout_c), .Q(i_4[3]));
    DFN1E1 \pd_pluse_data2[6]  (.D(pd_pluse_data[6]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[6]_net_1 ));
    DFN1E1 \pd_pluse_data3[2]  (.D(pd_pluse_data[2]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[2]_net_1 ));
    XA1A \pd_pluse_data2_RNIMASM[0]  (.A(\pd_pluse_data2[0]_net_1 ), 
        .B(count_5[0]), .C(\un1_count_3_i[0] ), .Y(\un1_count_NE_7[0] )
        );
    NOR3C \pd_pluse_data2_RNIC9791[12]  (.A(\un1_count_12_i[0] ), .B(
        \un1_count_9_i[0] ), .C(\un1_count_NE_7[0] ), .Y(
        \un1_count_NE_11[0] ));
    XNOR2 \pd_pluse_data1_RNIV2S6[14]  (.A(count_0[14]), .B(
        \pd_pluse_data1[14]_net_1 ), .Y(\i_reg10_14_i[0] ));
    NOR3A pd_pluse_data3_1_sqmuxa_0_a2_0 (.A(top_code_0_pd_pluse_load), 
        .B(pd_pluse_choice[3]), .C(pd_pluse_choice[2]), .Y(N_12));
    XNOR2 \pd_pluse_data1_RNINIR6[10]  (.A(count_0[10]), .B(
        \pd_pluse_data1[10]_net_1 ), .Y(\i_reg10_10_i[0] ));
    DFN1E1 \pd_pluse_data1[13]  (.D(pd_pluse_data[13]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[13]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3B pd_pluse_data2_1_sqmuxa_0_a2 (.A(pd_pluse_choice[1]), .B(
        N_12), .C(pd_pluse_choice[0]), .Y(pd_pluse_data2_1_sqmuxa));
    XA1A \pd_pluse_data1_RNI27TM[4]  (.A(\pd_pluse_data1[4]_net_1 ), 
        .B(count_5[4]), .C(\i_reg10_6_i[0] ), .Y(\i_reg10_NE_5[0] ));
    NOR3C \i_RNO_0[4]  (.A(\i_0_12[4] ), .B(\i_0_11[4] ), .C(
        \i_0_13[4] ), .Y(\i_0_15[4] ));
    DFN1E1 \pd_pluse_data2[7]  (.D(pd_pluse_data[7]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[7]_net_1 ));
    DFN1E1 \pd_pluse_data2[12]  (.D(pd_pluse_data[12]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[12]_net_1 ));
    DFN1E1 \pd_pluse_data1[3]  (.D(pd_pluse_data[3]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[3]_net_1 ));
    NOR2A \i_RNO[2]  (.A(net_27), .B(\i_reg10_NE[0] ), .Y(\i_RNO_2[2] )
        );
    NOR3C \pd_pluse_data2_RNIC9791[13]  (.A(\un1_count_1_0_i[0] ), .B(
        \un1_count_13_i[0] ), .C(\un1_count_NE_5[0] ), .Y(
        \un1_count_NE_10[0] ));
    NOR3C \i_RNO_12[4]  (.A(\un1_count_1_7_i_0[0] ), .B(
        \un1_count_1_5_i_0[0] ), .C(\i_0_4[4] ), .Y(\i_0_10[4] ));
    XA1A \pd_pluse_data2_RNI47TM[4]  (.A(\pd_pluse_data2[4]_net_1 ), 
        .B(count_5[4]), .C(\un1_count_6_i[0] ), .Y(\un1_count_NE_5[0] )
        );
    XNOR2 \pd_pluse_data2_RNI27S6[15]  (.A(count_0[15]), .B(
        \pd_pluse_data2[15]_net_1 ), .Y(\un1_count_15_i[0] ));
    DFN1E1 \pd_pluse_data2[9]  (.D(pd_pluse_data[9]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[9]_net_1 ));
    XNOR2 \pd_pluse_data1_RNINVEB[8]  (.A(count_0[8]), .B(
        \pd_pluse_data1[8]_net_1 ), .Y(\i_reg10_8_i[0] ));
    DFN1E1 \pd_pluse_data1[1]  (.D(pd_pluse_data[1]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[1]_net_1 ));
    NOR3C pd_pluse_data3_1_sqmuxa_0_a2 (.A(pd_pluse_choice[1]), .B(
        pd_pluse_choice[0]), .C(N_12), .Y(pd_pluse_data3_1_sqmuxa));
    DFN1E1 \pd_pluse_data3[8]  (.D(pd_pluse_data[8]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[8]_net_1 ));
    DFN1E1 \pd_pluse_data3[10]  (.D(pd_pluse_data[10]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[10]_net_1 ));
    XA1A \i_RNO_6[4]  (.A(\pd_pluse_data3[3]_net_1 ), .B(count_5[3]), 
        .C(\i_0_0[4] ), .Y(\i_0_8[4] ));
    OR2B \pd_pluse_data1_RNI8SOR4[11]  (.A(\i_reg10_NE_13[0] ), .B(
        \i_reg10_NE_12[0] ), .Y(\i_reg10_NE[0] ));
    DFN1E1 \pd_pluse_data3[13]  (.D(pd_pluse_data[13]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[13]_net_1 ));
    NOR3C \pd_pluse_data1_RNIGIEI2[13]  (.A(\i_reg10_NE_5[0] ), .B(
        \i_reg10_NE_4[0] ), .C(\i_reg10_NE_11[0] ), .Y(
        \i_reg10_NE_13[0] ));
    DFN1E1 \pd_pluse_data1[8]  (.D(pd_pluse_data[8]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[8]_net_1 ));
    NOR3C \pd_pluse_data2_RNI0AA92[2]  (.A(\un1_count_NE_3[0] ), .B(
        \un1_count_NE_2[0] ), .C(\un1_count_NE_8[0] ), .Y(
        \un1_count_NE_12[0] ));
    XA1A \pd_pluse_data1_RNICEAI[7]  (.A(\pd_pluse_data1[7]_net_1 ), 
        .B(count_2[7]), .C(\i_reg10_10_i[0] ), .Y(\i_reg10_NE_3[0] ));
    XNOR2 \pd_pluse_data1_RNIB7EB[2]  (.A(count_5[2]), .B(
        \pd_pluse_data1[2]_net_1 ), .Y(\i_reg10_2_i[0] ));
    DFN1E1 \pd_pluse_data3[5]  (.D(pd_pluse_data[5]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[5]_net_1 ));
    XA1A \pd_pluse_data2_RNIEEAI[7]  (.A(\pd_pluse_data2[7]_net_1 ), 
        .B(count_2[7]), .C(\un1_count_10_i[0] ), .Y(
        \un1_count_NE_3[0] ));
    XNOR2 \i_RNO_7[4]  (.A(count_5[4]), .B(\pd_pluse_data3[4]_net_1 ), 
        .Y(\un1_count_1_4_i_0[0] ));
    DFN1E1 \pd_pluse_data3[7]  (.D(pd_pluse_data[7]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[7]_net_1 ));
    NOR3C \pd_pluse_data2_RNIK0301[11]  (.A(\un1_count_8_i[0] ), .B(
        \un1_count_15_i[0] ), .C(\un1_count_NE_1[0] ), .Y(
        \un1_count_NE_8[0] ));
    XNOR2 \i_RNO_17[4]  (.A(count_2[7]), .B(\pd_pluse_data3[7]_net_1 ), 
        .Y(\un1_count_1_7_i_0[0] ));
    DFN1E1 \pd_pluse_data2[2]  (.D(pd_pluse_data[2]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[2]_net_1 ));
    DFN1E1 \pd_pluse_data1[9]  (.D(pd_pluse_data[9]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[9]_net_1 ));
    XNOR2 \pd_pluse_data2_RNIEBEB[3]  (.A(count_5[3]), .B(
        \pd_pluse_data2[3]_net_1 ), .Y(\un1_count_3_i[0] ));
    DFN1E1 \pd_pluse_data1[0]  (.D(pd_pluse_data[0]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[0]_net_1 ));
    XNOR2 \i_RNO_8[4]  (.A(count_5[1]), .B(\pd_pluse_data3[1]_net_1 ), 
        .Y(\un1_count_1_1_i_0[0] ));
    XNOR2 \i_RNO_18[4]  (.A(count_2[5]), .B(\pd_pluse_data3[5]_net_1 ), 
        .Y(\un1_count_1_5_i_0[0] ));
    NOR2B \i_RNO[0]  (.A(pulse_start_c), .B(net_27), .Y(\i_RNO_2[0] ));
    DFN1E1 \pd_pluse_data2[1]  (.D(pd_pluse_data[1]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[1]_net_1 ));
    DFN1E1 \pd_pluse_data2[0]  (.D(pd_pluse_data[0]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[0]_net_1 ));
    NOR3C \i_RNO_3[4]  (.A(\i_0_2[4] ), .B(\i_0_1[4] ), .C(\i_0_10[4] )
        , .Y(\i_0_13[4] ));
    DFN1 \i[0]  (.D(\i_RNO_2[0] ), .CLK(ddsclkout_c), .Q(i_5[0]));
    XNOR2 \pd_pluse_data2_RNIKNEB[6]  (.A(count_2[6]), .B(
        \pd_pluse_data2[6]_net_1 ), .Y(\un1_count_6_i[0] ));
    XNOR2 \pd_pluse_data1_RNIDBEB[3]  (.A(count_5[3]), .B(
        \pd_pluse_data1[3]_net_1 ), .Y(\i_reg10_3_i[0] ));
    XA1A \pd_pluse_data1_RNI62AI[13]  (.A(\pd_pluse_data1[13]_net_1 ), 
        .B(count_0[13]), .C(\i_reg10_1_i[0] ), .Y(\i_reg10_NE_4[0] ));
    DFN1E1 \pd_pluse_data1[14]  (.D(pd_pluse_data[14]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[14]_net_1 ));
    XNOR2 \i_RNO_5[4]  (.A(count_0[12]), .B(\pd_pluse_data3[12]_net_1 )
        , .Y(\un1_count_1_12_i_0[0] ));
    NOR3C \pd_pluse_data1_RNIO9A92[11]  (.A(\i_reg10_NE_1[0] ), .B(
        \i_reg10_NE_0[0] ), .C(\i_reg10_NE_9[0] ), .Y(
        \i_reg10_NE_12[0] ));
    DFN1E1 \pd_pluse_data2[8]  (.D(pd_pluse_data[8]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[8]_net_1 ));
    DFN1E1 \pd_pluse_data1[5]  (.D(pd_pluse_data[5]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[5]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1 \pd_pluse_data1[15]  (.D(pd_pluse_data[15]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[15]_net_1 ));
    XNOR2 \i_RNO_15[4]  (.A(count_5[2]), .B(\pd_pluse_data3[2]_net_1 ), 
        .Y(\un1_count_1_2_i_0[0] ));
    DFN1 \i[5]  (.D(\i_RNO_0[5] ), .CLK(ddsclkout_c), .Q(i_0[5]));
    XNOR2 \pd_pluse_data2_RNIIJEB[5]  (.A(count_2[5]), .B(
        \pd_pluse_data2[5]_net_1 ), .Y(\un1_count_5_i[0] ));
    DFN1E1 \pd_pluse_data1[11]  (.D(pd_pluse_data[11]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[11]_net_1 ));
    XNOR2 \pd_pluse_data1_RNIHJEB[5]  (.A(count_2[5]), .B(
        \pd_pluse_data1[5]_net_1 ), .Y(\i_reg10_5_i[0] ));
    XA1A \pd_pluse_data2_RNIUQSM[2]  (.A(\pd_pluse_data2[2]_net_1 ), 
        .B(count_5[2]), .C(\un1_count_5_i[0] ), .Y(\un1_count_NE_2[0] )
        );
    DFN1E1 \pd_pluse_data3[3]  (.D(pd_pluse_data[3]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[3]_net_1 ));
    NOR3C \pd_pluse_data1_RNI89791[12]  (.A(\i_reg10_12_i[0] ), .B(
        \i_reg10_9_i[0] ), .C(\i_reg10_NE_7[0] ), .Y(
        \i_reg10_NE_11[0] ));
    XNOR2 \pd_pluse_data2_RNIUUR6[13]  (.A(count_0[13]), .B(
        \pd_pluse_data2[13]_net_1 ), .Y(\un1_count_13_i[0] ));
    XNOR2 \pd_pluse_data2_RNIQ3FB[9]  (.A(count_0[9]), .B(
        \pd_pluse_data2[9]_net_1 ), .Y(\un1_count_9_i[0] ));
    XNOR2 \i_RNO_16[4]  (.A(count_0[11]), .B(
        \pd_pluse_data3[11]_net_1 ), .Y(\un1_count_1_11_i_0[0] ));
    XNOR2 \i_RNO_14[4]  (.A(count_0[9]), .B(\pd_pluse_data3[9]_net_1 ), 
        .Y(\un1_count_1_9_i_0[0] ));
    XNOR2 \pd_pluse_data2_RNI03S6[14]  (.A(count_0[14]), .B(
        \pd_pluse_data2[14]_net_1 ), .Y(\un1_count_14_i[0] ));
    XNOR2 \pd_pluse_data1_RNI93EB[1]  (.A(count_5[1]), .B(
        \pd_pluse_data1[1]_net_1 ), .Y(\i_reg10_1_i[0] ));
    DFN1E1 \pd_pluse_data3[14]  (.D(pd_pluse_data[14]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[14]_net_1 ));
    DFN1E1 \pd_pluse_data1[6]  (.D(pd_pluse_data[6]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[6]_net_1 ));
    XNOR2 \i_RNO_4[4]  (.A(count_5[0]), .B(\pd_pluse_data3[0]_net_1 ), 
        .Y(\un1_count_1_0_0_i_0[0] ));
    DFN1E1 \pd_pluse_data1[12]  (.D(pd_pluse_data[12]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[12]_net_1 ));
    XA1A \i_RNO_13[4]  (.A(\pd_pluse_data3[15]_net_1 ), .B(count_0[15])
        , .C(net_27), .Y(\i_0_0[4] ));
    XNOR2 \pd_pluse_data1_RNIJNEB[6]  (.A(count_2[6]), .B(
        \pd_pluse_data1[6]_net_1 ), .Y(\i_reg10_6_i[0] ));
    NOR3C \pd_pluse_data2_RNIOSOR4[12]  (.A(\un1_count_NE_11[0] ), .B(
        \un1_count_NE_10[0] ), .C(\un1_count_NE_12[0] ), .Y(
        \un1_count_i_i_0[0] ));
    DFN1E1 \pd_pluse_data2[4]  (.D(pd_pluse_data[4]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[4]_net_1 ));
    DFN1E1 \pd_pluse_data2[10]  (.D(pd_pluse_data[10]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[10]_net_1 ));
    DFN1E1 \pd_pluse_data3[15]  (.D(pd_pluse_data[15]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[15]_net_1 ));
    NOR3C \i_RNO_2[4]  (.A(\un1_count_1_4_i_0[0] ), .B(
        \un1_count_1_1_i_0[0] ), .C(\i_0_6[4] ), .Y(\i_0_11[4] ));
    DFN1E1 \pd_pluse_data2[3]  (.D(pd_pluse_data[3]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[3]_net_1 ));
    DFN1E1 \pd_pluse_data2[13]  (.D(pd_pluse_data[13]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[13]_net_1 ));
    DFN1E1 \pd_pluse_data3[11]  (.D(pd_pluse_data[11]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[11]_net_1 ));
    XA1A \i_RNO_10[4]  (.A(\pd_pluse_data3[14]_net_1 ), .B(count_0[14])
        , .C(\un1_count_1_2_i_0[0] ), .Y(\i_0_2[4] ));
    DFN1E1 \pd_pluse_data1[4]  (.D(pd_pluse_data[4]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[4]_net_1 ));
    XA1A \i_RNO_19[4]  (.A(\pd_pluse_data3[10]_net_1 ), .B(count_0[10])
        , .C(\un1_count_1_13_i_0[0] ), .Y(\i_0_4[4] ));
    XNOR2 \i_RNO_20[4]  (.A(count_0[13]), .B(
        \pd_pluse_data3[13]_net_1 ), .Y(\un1_count_1_13_i_0[0] ));
    DFN1E1 \pd_pluse_data3[12]  (.D(pd_pluse_data[12]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[12]_net_1 ));
    XNOR2 \pd_pluse_data2_RNIA3EB[1]  (.A(count_5[1]), .B(
        \pd_pluse_data2[1]_net_1 ), .Y(\un1_count_1_0_i[0] ));
    NOR3C \i_RNO_1[4]  (.A(\un1_count_1_0_0_i_0[0] ), .B(
        \un1_count_1_12_i_0[0] ), .C(\i_0_8[4] ), .Y(\i_0_12[4] ));
    XA1A \pd_pluse_data1_RNIKASM[0]  (.A(\pd_pluse_data1[0]_net_1 ), 
        .B(count_5[0]), .C(\i_reg10_3_i[0] ), .Y(\i_reg10_NE_7[0] ));
    DFN1 \i[4]  (.D(\i_RNO_0[4]_net_1 ), .CLK(ddsclkout_c), .Q(i_0[4]));
    XNOR2 \pd_pluse_data2_RNIOIR6[10]  (.A(count_0[10]), .B(
        \pd_pluse_data2[10]_net_1 ), .Y(\un1_count_10_i[0] ));
    XNOR2 \pd_pluse_data1_RNIP3FB[9]  (.A(count_0[9]), .B(
        \pd_pluse_data1[9]_net_1 ), .Y(\i_reg10_9_i[0] ));
    DFN1E1 \pd_pluse_data2[5]  (.D(pd_pluse_data[5]), .CLK(GLA), .E(
        pd_pluse_data2_1_sqmuxa), .Q(\pd_pluse_data2[5]_net_1 ));
    DFN1E1 \pd_pluse_data1[2]  (.D(pd_pluse_data[2]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[2]_net_1 ));
    XA1A \i_RNO_9[4]  (.A(\pd_pluse_data3[6]_net_1 ), .B(count_2[6]), 
        .C(\un1_count_1_9_i_0[0] ), .Y(\i_0_6[4] ));
    NOR2B \i_RNO[5]  (.A(net_27), .B(bri_dump_sw_0_tetw_pluse), .Y(
        \i_RNO_0[5] ));
    DFN1E1 \pd_pluse_data3[4]  (.D(pd_pluse_data[4]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[4]_net_1 ));
    DFN1E1 \pd_pluse_data3[1]  (.D(pd_pluse_data[1]), .CLK(GLA), .E(
        pd_pluse_data3_1_sqmuxa), .Q(\pd_pluse_data3[1]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1E1 \pd_pluse_data1[7]  (.D(pd_pluse_data[7]), .CLK(GLA), .E(
        pd_pluse_data1_0_sqmuxa), .Q(\pd_pluse_data1[7]_net_1 ));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module pd_pluse_state(
       i_5,
       i_0,
       i_4,
       pd_pulse_en_c,
       ddsclkout_c,
       pd_pluse_state_0_stateover,
       net_27
    );
input  [0:0] i_5;
input  [5:4] i_0;
input  [3:1] i_4;
output pd_pulse_en_c;
input  ddsclkout_c;
output pd_pluse_state_0_stateover;
input  net_27;

    wire en1_0_i_0, N_166, cs_1, \cs_srsts_0_i_a5_1[12] , 
        \cs[11]_net_1 , \cs[12]_net_1 , \cs_srsts_0_i_a5_0[12] , 
        \cs[4]_net_1 , \cs[7]_net_1 , N_195, en1_RNO_net_1, N_184, 
        N_183, \cs_RNO_0[9]_net_1 , N_178, N_177, \cs_RNO_1[8] , 
        \cs_i[0]_net_1 , \cs_RNO_1[7] , en2, \cs_RNO_3[3] , N_175, 
        N_174, \cs[9]_net_1 , \cs[2]_net_1 , \cs_RNO[10]_net_1 , N_180, 
        N_179, \cs_RNO_2[6] , N_185, N_186, \cs[3]_net_1 , 
        \cs_RNO_2[1] , \cs[8]_net_1 , \cs_RNO_1[2] , N_168, N_167, 
        \cs_RNO_3[5] , N_170, \cs[5]_net_1 , \cs_RNO_1[12] , 
        \cs[1]_net_1 , en_RNO_net_1, en1_net_1, stateover_RNO_1, 
        \cs_RNO_2[4] , \cs_RNO_1[11] , \cs[10]_net_1 , GND, VCC, GND_0, 
        VCC_0;
    
    NOR3A \cs_RNO[10]  (.A(cs_1), .B(N_180), .C(N_179), .Y(
        \cs_RNO[10]_net_1 ));
    DFN1 \cs[6]  (.D(\cs_RNO_2[6] ), .CLK(ddsclkout_c), .Q(en2));
    NOR3C \cs_RNO[11]  (.A(cs_1), .B(i_4[3]), .C(\cs[10]_net_1 ), .Y(
        \cs_RNO_1[11] ));
    AOI1 \cs_RNO_1[3]  (.A(i_4[2]), .B(\cs[2]_net_1 ), .C(
        \cs[3]_net_1 ), .Y(N_174));
    DFN1 \cs[12]  (.D(\cs_RNO_1[12] ), .CLK(ddsclkout_c), .Q(
        \cs[12]_net_1 ));
    NOR2 en1_RNO_1 (.A(i_4[2]), .B(N_166), .Y(N_183));
    VCC VCC_i (.Y(VCC));
    OR2 \cs_RNI8N7A[3]  (.A(\cs[10]_net_1 ), .B(\cs[3]_net_1 ), .Y(
        N_166));
    DFN1 \cs[3]  (.D(\cs_RNO_3[3] ), .CLK(ddsclkout_c), .Q(
        \cs[3]_net_1 ));
    NOR3C \cs_RNO[7]  (.A(en2), .B(i_0[4]), .C(cs_1), .Y(\cs_RNO_1[7] )
        );
    NOR2B \cs_RNO[1]  (.A(\cs[8]_net_1 ), .B(cs_1), .Y(\cs_RNO_2[1] ));
    NOR3A \cs_RNO[9]  (.A(cs_1), .B(N_178), .C(N_177), .Y(
        \cs_RNO_0[9]_net_1 ));
    DFN1 \cs[5]  (.D(\cs_RNO_3[5] ), .CLK(ddsclkout_c), .Q(
        \cs[5]_net_1 ));
    OA1 en_RNO (.A(en1_net_1), .B(en2), .C(cs_1), .Y(en_RNO_net_1));
    NOR2A \cs_RNO_0[3]  (.A(i_4[3]), .B(\cs[2]_net_1 ), .Y(N_175));
    NOR3B \cs_RNO[8]  (.A(i_0[5]), .B(cs_1), .C(\cs_i[0]_net_1 ), .Y(
        \cs_RNO_1[8] ));
    OR2 \cs_RNIVTE9[4]  (.A(\cs[4]_net_1 ), .B(\cs[7]_net_1 ), .Y(
        \cs_srsts_0_i_a5_0[12] ));
    DFN1 \cs[11]  (.D(\cs_RNO_1[11] ), .CLK(ddsclkout_c), .Q(
        \cs[11]_net_1 ));
    OA1A \cs_RNO_1[9]  (.A(\cs[9]_net_1 ), .B(i_4[2]), .C(
        \cs_i[0]_net_1 ), .Y(N_177));
    DFN1 \cs[2]  (.D(\cs_RNO_1[2] ), .CLK(ddsclkout_c), .Q(
        \cs[2]_net_1 ));
    DFN1 en1 (.D(en1_RNO_net_1), .CLK(ddsclkout_c), .Q(en1_net_1));
    NOR3 en1_RNO (.A(N_184), .B(N_183), .C(en1_0_i_0), .Y(
        en1_RNO_net_1));
    DFN1 en (.D(en_RNO_net_1), .CLK(ddsclkout_c), .Q(pd_pulse_en_c));
    NOR2A \cs_RNO[12]  (.A(cs_1), .B(N_195), .Y(\cs_RNO_1[12] ));
    GND GND_i (.Y(GND));
    NOR2 \cs_RNO_0[10]  (.A(i_4[2]), .B(\cs[10]_net_1 ), .Y(N_180));
    NOR2B un1_state_initial_0_o5 (.A(i_5[0]), .B(net_27), .Y(cs_1));
    DFN1 \cs_i[0]  (.D(cs_1), .CLK(ddsclkout_c), .Q(\cs_i[0]_net_1 ));
    DFN1 stateover (.D(stateover_RNO_1), .CLK(ddsclkout_c), .Q(
        pd_pluse_state_0_stateover));
    AO1C \cs_RNIR6A9[1]  (.A(\cs[1]_net_1 ), .B(i_4[2]), .C(cs_1), .Y(
        N_167));
    DFN1 \cs[10]  (.D(\cs_RNO[10]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[10]_net_1 ));
    NOR2 \cs_RNO_0[6]  (.A(i_4[2]), .B(en2), .Y(N_185));
    OA1B \cs_RNO[2]  (.A(N_168), .B(\cs[2]_net_1 ), .C(N_167), .Y(
        \cs_RNO_1[2] ));
    OA1C \cs_RNO_1[10]  (.A(\cs[10]_net_1 ), .B(i_4[3]), .C(
        \cs[9]_net_1 ), .Y(N_179));
    NOR2A \cs_RNO_0[2]  (.A(\cs[1]_net_1 ), .B(i_4[1]), .Y(N_168));
    OR2 \cs_RNIPS0B[11]  (.A(\cs[11]_net_1 ), .B(\cs[12]_net_1 ), .Y(
        \cs_srsts_0_i_a5_1[12] ));
    AO1B stateover_RNO (.A(pd_pluse_state_0_stateover), .B(N_195), .C(
        cs_1), .Y(stateover_RNO_1));
    NOR3 en1_RNO_0 (.A(\cs[9]_net_1 ), .B(\cs[2]_net_1 ), .C(N_166), 
        .Y(N_184));
    NOR3C \cs_RNO[4]  (.A(cs_1), .B(i_4[3]), .C(\cs[3]_net_1 ), .Y(
        \cs_RNO_2[4] ));
    DFN1 \cs[9]  (.D(\cs_RNO_0[9]_net_1 ), .CLK(ddsclkout_c), .Q(
        \cs[9]_net_1 ));
    NOR2B \cs_RNO_0[5]  (.A(i_4[1]), .B(\cs[1]_net_1 ), .Y(N_170));
    DFN1 \cs[8]  (.D(\cs_RNO_1[8] ), .CLK(ddsclkout_c), .Q(
        \cs[8]_net_1 ));
    OA1C \cs_RNO_1[6]  (.A(en2), .B(i_0[4]), .C(\cs[5]_net_1 ), .Y(
        N_186));
    NOR3A \cs_RNO[6]  (.A(cs_1), .B(N_185), .C(N_186), .Y(
        \cs_RNO_2[6] ));
    NOR2 \cs_RNIOQFK[4]  (.A(\cs_srsts_0_i_a5_1[12] ), .B(
        \cs_srsts_0_i_a5_0[12] ), .Y(N_195));
    NOR3A \cs_RNO[3]  (.A(cs_1), .B(N_175), .C(N_174), .Y(
        \cs_RNO_3[3] ));
    DFN1 \cs[1]  (.D(\cs_RNO_2[1] ), .CLK(ddsclkout_c), .Q(
        \cs[1]_net_1 ));
    OA1B \cs_RNO[5]  (.A(N_170), .B(\cs[5]_net_1 ), .C(N_167), .Y(
        \cs_RNO_3[5] ));
    DFN1 \cs[4]  (.D(\cs_RNO_2[4] ), .CLK(ddsclkout_c), .Q(
        \cs[4]_net_1 ));
    DFN1 \cs[7]  (.D(\cs_RNO_1[7] ), .CLK(ddsclkout_c), .Q(
        \cs[7]_net_1 ));
    AO1B en1_RNO_2 (.A(i_4[3]), .B(N_166), .C(cs_1), .Y(en1_0_i_0));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    NOR2A \cs_RNO_0[9]  (.A(i_0[5]), .B(\cs[9]_net_1 ), .Y(N_178));
    
endmodule


module pd_pluse_inc(
       count_2,
       count_5,
       count_0,
       count1
    );
input  [7:5] count_2;
input  [4:0] count_5;
input  [15:8] count_0;
output [15:1] count1;

    wire Rcout_8_net, Rcout_5_net, inc_2_net, Rcout_6_net, inc_5_net, 
        Rcout_13_net, inc_17_net, inc_16_net, Rcout_4_net, inc_20_net, 
        Rcout_12_net, Rcout_14_net, Rcout_10_net, inc_12_net, 
        inc_10_net, Rcout_11_net, inc_14_net, Rcout_9_net, incb_2_net, 
        inc_22_net, incb_5_net, Rcout_15_net, inc_1_net, inc_8_net, 
        Rcout_7_net, GND, VCC, GND_0, VCC_0;
    
    AND3 AND2b_9_inst (.A(count_5[0]), .B(count_5[1]), .C(count_5[2]), 
        .Y(incb_2_net));
    AND3 FND2_9_inst (.A(inc_12_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_10_net));
    AND2 AND2_4_inst (.A(inc_2_net), .B(count_5[3]), .Y(Rcout_4_net));
    AND3 AND2_15_inst (.A(inc_16_net), .B(inc_17_net), .C(inc_20_net), 
        .Y(Rcout_14_net));
    AND3 AND2_1_12_inst (.A(incb_2_net), .B(incb_5_net), .C(inc_10_net)
        , .Y(inc_17_net));
    AND2 AND2_13_inst (.A(inc_17_net), .B(inc_16_net), .Y(Rcout_12_net)
        );
    AND3 AND2_12_inst (.A(count_0[9]), .B(count_0[10]), .C(count_0[11])
        , .Y(inc_16_net));
    VCC VCC_i (.Y(VCC));
    AND3 AND2_1_7_inst (.A(inc_2_net), .B(inc_5_net), .C(count_2[6]), 
        .Y(Rcout_7_net));
    XOR2 HOR2_10_inst (.A(Rcout_13_net), .B(count_0[13]), .Y(
        count1[13]));
    AND3 AND2_1_8_inst (.A(inc_2_net), .B(inc_5_net), .C(inc_8_net), 
        .Y(Rcout_8_net));
    XOR2 XOR2_4_inst (.A(Rcout_5_net), .B(count_2[5]), .Y(count1[5]));
    AND2 AND2_7_inst (.A(inc_2_net), .B(inc_5_net), .Y(Rcout_6_net));
    AND2 AND2_14_inst (.A(count_0[12]), .B(count_0[13]), .Y(inc_20_net)
        );
    AND3 TND2_15_inst (.A(inc_16_net), .B(inc_17_net), .C(inc_22_net), 
        .Y(Rcout_15_net));
    XOR2 XOR2_3_inst (.A(Rcout_4_net), .B(count_5[4]), .Y(count1[4]));
    AND2 FND2_8_inst (.A(incb_2_net), .B(count_0[9]), .Y(inc_12_net));
    XOR2 XOR2_7_inst (.A(Rcout_9_net), .B(count_0[9]), .Y(count1[9]));
    XOR2 UXOR2_12_inst (.A(Rcout_15_net), .B(count_0[15]), .Y(
        count1[15]));
    AND3 AND2_9_inst (.A(count_2[6]), .B(count_2[7]), .C(count_0[8]), 
        .Y(inc_10_net));
    GND GND_i (.Y(GND));
    AND3 AND2_11_inst (.A(inc_14_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_11_net));
    XOR2 XOR2_6_inst (.A(Rcout_8_net), .B(count_0[8]), .Y(count1[8]));
    XOR2 XOR2_1_5_inst (.A(Rcout_7_net), .B(count_2[7]), .Y(count1[7]));
    AND3 TAND2_15_inst (.A(count_0[12]), .B(count_0[13]), .C(
        count_0[14]), .Y(inc_22_net));
    AND3 AND2_3_inst (.A(count_5[0]), .B(count_5[1]), .C(count_5[2]), 
        .Y(inc_2_net));
    AND3 fAND2_8_inst (.A(incb_2_net), .B(inc_5_net), .C(inc_10_net), 
        .Y(Rcout_9_net));
    AND3 AND2_6_inst (.A(count_5[3]), .B(count_5[4]), .C(count_2[5]), 
        .Y(inc_5_net));
    AND3 AND2b_12_inst (.A(count_5[3]), .B(count_5[4]), .C(count_2[5]), 
        .Y(incb_5_net));
    XOR2 XOR2_2_1_inst (.A(inc_1_net), .B(count_5[2]), .Y(count1[2]));
    XOR2 XOR2_1_inst (.A(count_5[0]), .B(count_5[1]), .Y(count1[1]));
    XOR2 XOR2_9_inst (.A(Rcout_11_net), .B(count_0[11]), .Y(count1[11])
        );
    XOR2 XOR2_2_inst (.A(inc_2_net), .B(count_5[3]), .Y(count1[3]));
    AND2 AND2_8_inst (.A(count_2[6]), .B(count_2[7]), .Y(inc_8_net));
    AND3 HND2_13_inst (.A(inc_17_net), .B(inc_16_net), .C(count_0[12]), 
        .Y(Rcout_13_net));
    XOR2 POR2_9_inst (.A(Rcout_12_net), .B(count_0[12]), .Y(count1[12])
        );
    XOR2 XOR2_5_inst (.A(Rcout_6_net), .B(count_2[6]), .Y(count1[6]));
    AND2 AND2_2_inst (.A(count_5[0]), .B(count_5[1]), .Y(inc_1_net));
    AND3 AND2_5_inst (.A(inc_2_net), .B(count_5[3]), .C(count_5[4]), 
        .Y(Rcout_5_net));
    XOR2 FOR2_8_inst (.A(Rcout_10_net), .B(count_0[10]), .Y(count1[10])
        );
    XOR2 XOR2_11_inst (.A(Rcout_14_net), .B(count_0[14]), .Y(
        count1[14]));
    AND3 AND2_10_inst (.A(incb_2_net), .B(count_0[9]), .C(count_0[10]), 
        .Y(inc_14_net));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module pd_pluse_timer(
       count_0,
       count_2,
       count_5,
       net_27,
       ddsclkout_c,
       pulse_start_c,
       pd_pluse_state_0_stateover
    );
output [15:8] count_0;
output [7:5] count_2;
output [4:0] count_5;
input  net_27;
input  ddsclkout_c;
input  pulse_start_c;
input  pd_pluse_state_0_stateover;

    wire \count_3[0] , \count_3[1] , \count1[1] , \count_3[2] , 
        \count1[2] , \count_3[3] , \count1[3] , \count_3[4] , 
        \count1[4] , \count_3[5] , \count1[5] , \count_3[6] , 
        \count1[6] , \count_3[7] , \count1[7] , \count_3[8] , 
        \count1[8] , \count_3[9] , \count1[9] , \count_3[10] , 
        \count1[10] , \count_3[11] , \count1[11] , \count_3[12] , 
        \count1[12] , \count_3[13] , \count1[13] , \count_3[14] , 
        \count1[14] , \count_3[15] , \count1[15] , GND, VCC, GND_0, 
        VCC_0;
    
    DFN1C0 \count[5]  (.D(\count_3[5] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_2[5]));
    DFN1C0 \count[1]  (.D(\count_3[1] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_5[1]));
    DFN1C0 \count[10]  (.D(\count_3[10] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[10]));
    DFN1C0 \count[0]  (.D(\count_3[0] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_5[0]));
    DFN1C0 \count[14]  (.D(\count_3[14] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[14]));
    NOR3C \count_RNO[7]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[7] ), .Y(\count_3[7] ));
    NOR3C \count_RNO[15]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[15] ), .Y(\count_3[15] ));
    NOR3C \count_RNO[2]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[2] ), .Y(\count_3[2] ));
    NOR3C \count_RNO[9]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[9] ), .Y(\count_3[9] ));
    VCC VCC_i (.Y(VCC));
    NOR3C \count_RNO[4]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[4] ), .Y(\count_3[4] ));
    DFN1C0 \count[8]  (.D(\count_3[8] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[8]));
    NOR3C \count_RNO[10]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[10] ), .Y(\count_3[10] ));
    DFN1C0 \count[15]  (.D(\count_3[15] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[15]));
    NOR3C \count_RNO[3]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[3] ), .Y(\count_3[3] ));
    DFN1C0 \count[11]  (.D(\count_3[11] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[11]));
    NOR3C \count_RNO[8]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[8] ), .Y(\count_3[8] ));
    DFN1C0 \count[13]  (.D(\count_3[13] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[13]));
    NOR3C \count_RNO[5]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[5] ), .Y(\count_3[5] ));
    NOR3C \count_RNO[1]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[1] ), .Y(\count_3[1] ));
    NOR3C \count_RNO[11]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[11] ), .Y(\count_3[11] ));
    DFN1C0 \count[2]  (.D(\count_3[2] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_5[2]));
    pd_pluse_inc pd_pluse_inc_0 (.count_2({count_2[7], count_2[6], 
        count_2[5]}), .count_5({count_5[4], count_5[3], count_5[2], 
        count_5[1], count_5[0]}), .count_0({count_0[15], count_0[14], 
        count_0[13], count_0[12], count_0[11], count_0[10], count_0[9], 
        count_0[8]}), .count1({\count1[15] , \count1[14] , 
        \count1[13] , \count1[12] , \count1[11] , \count1[10] , 
        \count1[9] , \count1[8] , \count1[7] , \count1[6] , 
        \count1[5] , \count1[4] , \count1[3] , \count1[2] , 
        \count1[1] }));
    GND GND_i (.Y(GND));
    DFN1C0 \count[9]  (.D(\count_3[9] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[9]));
    NOR3C \count_RNO[6]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[6] ), .Y(\count_3[6] ));
    NOR3C \count_RNO[12]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[12] ), .Y(\count_3[12] ));
    NOR3B \count_RNO[0]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(count_5[0]), .Y(\count_3[0] ));
    DFN1C0 \count[6]  (.D(\count_3[6] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_2[6]));
    DFN1C0 \count[3]  (.D(\count_3[3] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_5[3]));
    NOR3C \count_RNO[14]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[14] ), .Y(\count_3[14] ));
    NOR3C \count_RNO[13]  (.A(pd_pluse_state_0_stateover), .B(
        pulse_start_c), .C(\count1[13] ), .Y(\count_3[13] ));
    DFN1C0 \count[4]  (.D(\count_3[4] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_5[4]));
    DFN1C0 \count[12]  (.D(\count_3[12] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_0[12]));
    DFN1C0 \count[7]  (.D(\count_3[7] ), .CLK(ddsclkout_c), .CLR(
        net_27), .Q(count_2[7]));
    VCC VCC_i_0 (.Y(VCC_0));
    GND GND_i_0 (.Y(GND_0));
    
endmodule


module pd_pluse_top(
       i_4_0,
       pd_pluse_choice,
       i_0_0,
       pd_pluse_data,
       pd_pulse_en_c,
       net_27,
       top_code_0_pd_pluse_load,
       pulse_start_c,
       net_51,
       bri_dump_sw_0_tetw_pluse,
       GLA,
       ddsclkout_c
    );
input  i_4_0;
input  [3:0] pd_pluse_choice;
output [1:1] i_0_0;
input  [15:0] pd_pluse_data;
output pd_pulse_en_c;
input  net_27;
input  top_code_0_pd_pluse_load;
input  pulse_start_c;
input  net_51;
input  bri_dump_sw_0_tetw_pluse;
input  GLA;
input  ddsclkout_c;

    wire \i_0[4] , \i_0[5] , \i_4[2] , \i_4[3] , \i_5[0] , 
        \count_0[8] , \count_0[9] , \count_0[10] , \count_0[11] , 
        \count_0[12] , \count_0[13] , \count_0[14] , \count_0[15] , 
        \count_2[5] , \count_2[6] , \count_2[7] , \count_5[0] , 
        \count_5[1] , \count_5[2] , \count_5[3] , \count_5[4] , 
        pd_pluse_state_0_stateover, GND, VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    pd_pluse_coder pd_pluse_coder_0 (.i_0({\i_0[5] , \i_0[4] }), .i_4({
        \i_4[3] , \i_4[2] }), .i_5({\i_5[0] }), .pd_pluse_data({
        pd_pluse_data[15], pd_pluse_data[14], pd_pluse_data[13], 
        pd_pluse_data[12], pd_pluse_data[11], pd_pluse_data[10], 
        pd_pluse_data[9], pd_pluse_data[8], pd_pluse_data[7], 
        pd_pluse_data[6], pd_pluse_data[5], pd_pluse_data[4], 
        pd_pluse_data[3], pd_pluse_data[2], pd_pluse_data[1], 
        pd_pluse_data[0]}), .i_0_0_0(i_0_0[1]), .pd_pluse_choice({
        pd_pluse_choice[3], pd_pluse_choice[2], pd_pluse_choice[1], 
        pd_pluse_choice[0]}), .count_0({\count_0[15] , \count_0[14] , 
        \count_0[13] , \count_0[12] , \count_0[11] , \count_0[10] , 
        \count_0[9] , \count_0[8] }), .count_2({\count_2[7] , 
        \count_2[6] , \count_2[5] }), .count_5({\count_5[4] , 
        \count_5[3] , \count_5[2] , \count_5[1] , \count_5[0] }), 
        .ddsclkout_c(ddsclkout_c), .GLA(GLA), 
        .bri_dump_sw_0_tetw_pluse(bri_dump_sw_0_tetw_pluse), .net_51(
        net_51), .pulse_start_c(pulse_start_c), 
        .top_code_0_pd_pluse_load(top_code_0_pd_pluse_load), .net_27(
        net_27));
    pd_pluse_state pd_pluse_state_0 (.i_5({\i_5[0] }), .i_0({\i_0[5] , 
        \i_0[4] }), .i_4({\i_4[3] , \i_4[2] , i_4_0}), .pd_pulse_en_c(
        pd_pulse_en_c), .ddsclkout_c(ddsclkout_c), 
        .pd_pluse_state_0_stateover(pd_pluse_state_0_stateover), 
        .net_27(net_27));
    GND GND_i_0 (.Y(GND_0));
    pd_pluse_timer pd_pluse_timer_0 (.count_0({\count_0[15] , 
        \count_0[14] , \count_0[13] , \count_0[12] , \count_0[11] , 
        \count_0[10] , \count_0[9] , \count_0[8] }), .count_2({
        \count_2[7] , \count_2[6] , \count_2[5] }), .count_5({
        \count_5[4] , \count_5[3] , \count_5[2] , \count_5[1] , 
        \count_5[0] }), .net_27(net_27), .ddsclkout_c(ddsclkout_c), 
        .pulse_start_c(pulse_start_c), .pd_pluse_state_0_stateover(
        pd_pluse_state_0_stateover));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_1(
       i_5,
       i_6,
       GLA,
       off_on_state_0_state_over,
       DUMP_ON_0_dump_on,
       OR2_2_Y
    );
input  [1:1] i_5;
input  [0:0] i_6;
input  GLA;
output off_on_state_0_state_over;
output DUMP_ON_0_dump_on;
input  OR2_2_Y;

    wire N_14, N_13, \cs_nsss[0] , N_42, \cs_nsss[1] , \cs_ns[1] , 
        \cs[1]_net_1 , GND, VCC, GND_0, VCC_0;
    
    OR2B state_over_RNO_0 (.A(off_on_state_0_state_over), .B(N_42), .Y(
        N_13));
    DFN1 state_over (.D(N_14), .CLK(GLA), .Q(off_on_state_0_state_over)
        );
    DFN1 \cs[0]  (.D(\cs_nsss[0] ), .CLK(GLA), .Q(DUMP_ON_0_dump_on));
    NOR3C \cs_RNO[0]  (.A(N_42), .B(OR2_2_Y), .C(i_6[0]), .Y(
        \cs_nsss[0] ));
    AOI1 \cs_RNISLRA[1]  (.A(DUMP_ON_0_dump_on), .B(i_5[1]), .C(
        \cs[1]_net_1 ), .Y(N_42));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 \cs[1]  (.D(\cs_nsss[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3C \cs_RNO[1]  (.A(\cs_ns[1] ), .B(OR2_2_Y), .C(i_6[0]), .Y(
        \cs_nsss[1] ));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    MX2 \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_5[1]), .S(
        DUMP_ON_0_dump_on), .Y(\cs_ns[1] ));
    OR3C state_over_RNO (.A(N_13), .B(i_6[0]), .C(OR2_2_Y), .Y(N_14));
    
endmodule


module off_on_coder_1(
       i_5,
       i_6,
       count_6,
       GLA,
       OR2_1_Y,
       OR2_2_Y
    );
output [1:1] i_5;
output [0:0] i_6;
input  [4:0] count_6;
input  GLA;
input  OR2_1_Y;
input  OR2_2_Y;

    wire \i_0_1[1] , \i_RNO_2[1] , N_17, \i_RNO_3[0] , GND, VCC, GND_0, 
        VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \i_RNO_1[1]  (.A(count_6[1]), .B(count_6[0]), .Y(N_17));
    DFN1 \i[1]  (.D(\i_RNO_2[1] ), .CLK(GLA), .Q(i_5[1]));
    GND GND_i_0 (.Y(GND_0));
    NOR3C \i_RNO[1]  (.A(\i_0_1[1] ), .B(N_17), .C(OR2_2_Y), .Y(
        \i_RNO_2[1] ));
    VCC VCC_i (.Y(VCC));
    NOR3B \i_RNO_0[1]  (.A(count_6[2]), .B(count_6[4]), .C(count_6[3]), 
        .Y(\i_0_1[1] ));
    NOR2B \i_RNO[0]  (.A(OR2_2_Y), .B(OR2_1_Y), .Y(\i_RNO_3[0] ));
    DFN1 \i[0]  (.D(\i_RNO_3[0] ), .CLK(GLA), .Q(i_6[0]));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_1(
       count_6,
       GLA,
       OR2_2_Y,
       off_on_state_0_state_over,
       OR2_1_Y
    );
output [4:0] count_6;
input  GLA;
input  OR2_2_Y;
input  off_on_state_0_state_over;
input  OR2_1_Y;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_15_i, GND, VCC, GND_0, VCC_0;
    
    NOR2B \count_RNILBUF[1]  (.A(count_6[1]), .B(count_6[0]), .Y(N_12));
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_6[0]), .B(count_6[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_6[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_6[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count_6[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    VCC VCC_i (.Y(VCC));
    NOR2B \count_RNIHHTN[2]  (.A(count_6[2]), .B(N_12), .Y(N_13));
    GND GND_i (.Y(GND));
    AX1E \count_RNO_0[4]  (.A(N_13), .B(count_6[3]), .C(count_6[4]), 
        .Y(N_15_i));
    XA1B \count_RNO[2]  (.A(N_12), .B(count_6[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(OR2_1_Y), .B(off_on_state_0_state_over), 
        .C(OR2_2_Y), .Y(count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \count_RNO[4]  (.A(count_0_sqmuxa_net_1), .B(N_15_i), .Y(N_11)
        );
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_6[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_6[4]));
    NOR2 \count_RNO[0]  (.A(count_6[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_6[2]));
    
endmodule


module DUMP_ON(
       OR2_1_Y,
       OR2_2_Y,
       DUMP_ON_0_dump_on,
       GLA
    );
input  OR2_1_Y;
input  OR2_2_Y;
output DUMP_ON_0_dump_on;
input  GLA;

    wire \i_5[1] , \i_6[0] , off_on_state_0_state_over, \count_6[0] , 
        \count_6[1] , \count_6[2] , \count_6[3] , \count_6[4] , GND, 
        VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1_1 
        off_on_state_0 (.i_5({\i_5[1] }), .i_6({\i_6[0] }), .GLA(GLA), 
        .off_on_state_0_state_over(off_on_state_0_state_over), 
        .DUMP_ON_0_dump_on(DUMP_ON_0_dump_on), .OR2_2_Y(OR2_2_Y));
    off_on_coder_1 off_on_coder_0 (.i_5({\i_5[1] }), .i_6({\i_6[0] }), 
        .count_6({\count_6[4] , \count_6[3] , \count_6[2] , 
        \count_6[1] , \count_6[0] }), .GLA(GLA), .OR2_1_Y(OR2_1_Y), 
        .OR2_2_Y(OR2_2_Y));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0_1 
        off_on_timer_0 (.count_6({\count_6[4] , \count_6[3] , 
        \count_6[2] , \count_6[1] , \count_6[0] }), .GLA(GLA), 
        .OR2_2_Y(OR2_2_Y), .off_on_state_0_state_over(
        off_on_state_0_state_over), .OR2_1_Y(OR2_1_Y));
    GND GND_i (.Y(GND));
    
endmodule


module nsctrl_choice(
       nsctrl_choice_0_dumpoff_ctr,
       nsctrl_choice_0_dumpon_ctr,
       nsctrl_choice_0_dumponoff_rst,
       nsctrl_choice_0_intertodsp,
       nsctrl_choice_0_rt_sw,
       nsctrl_choice_0_soft_d,
       GLA,
       nsctrl_choice_0_sw_acq2,
       noisestate_0_sw_acq2,
       scanstate_0_sw_acq2,
       top_code_0_n_s_ctrl,
       noisestate_0_rt_sw,
       scanstate_0_rt_sw,
       noisestate_0_dumpon_ctr,
       scanstate_0_dds_conf,
       top_code_0_n_s_ctrl_1,
       noisestate_0_soft_d,
       scanstate_0_soft_d,
       noisestate_0_state_over_n,
       scanstate_0_state_over_n,
       top_code_0_noise_rst_0,
       net_33_0,
       top_code_0_n_s_ctrl_0,
       noisestate_0_dumpoff_ctr,
       scanstate_0_dumpoff_ctr,
       net_27
    );
output nsctrl_choice_0_dumpoff_ctr;
output nsctrl_choice_0_dumpon_ctr;
output nsctrl_choice_0_dumponoff_rst;
output nsctrl_choice_0_intertodsp;
output nsctrl_choice_0_rt_sw;
output nsctrl_choice_0_soft_d;
input  GLA;
output nsctrl_choice_0_sw_acq2;
input  noisestate_0_sw_acq2;
input  scanstate_0_sw_acq2;
input  top_code_0_n_s_ctrl;
input  noisestate_0_rt_sw;
input  scanstate_0_rt_sw;
input  noisestate_0_dumpon_ctr;
input  scanstate_0_dds_conf;
input  top_code_0_n_s_ctrl_1;
input  noisestate_0_soft_d;
input  scanstate_0_soft_d;
input  noisestate_0_state_over_n;
input  scanstate_0_state_over_n;
input  top_code_0_noise_rst_0;
input  net_33_0;
input  top_code_0_n_s_ctrl_0;
input  noisestate_0_dumpoff_ctr;
input  scanstate_0_dumpoff_ctr;
input  net_27;

    wire intertodsp_RNO_net_1, intertodsp_5, dumponoff_rst_RNO_net_1, 
        dumponoff_rst_5, dumpoff_ctr_RNO_net_1, dumpoff_ctr_5, 
        soft_d_5, dumpon_ctr_5, dumpon_ctr_RNO_net_1, soft_d_RNO_net_1, 
        rt_sw_5, rt_sw_RNO_net_1, sw_acq2_5, sw_acq2_RNO_net_1, GND, 
        VCC, GND_0, VCC_0;
    
    MX2C sw_acq2_RNO_0 (.A(scanstate_0_sw_acq2), .B(
        noisestate_0_sw_acq2), .S(top_code_0_n_s_ctrl), .Y(sw_acq2_5));
    DFN1 rt_sw (.D(rt_sw_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_rt_sw));
    NOR2A dumpon_ctr_RNO (.A(net_27), .B(dumpon_ctr_5), .Y(
        dumpon_ctr_RNO_net_1));
    MX2C rt_sw_RNO_0 (.A(scanstate_0_rt_sw), .B(noisestate_0_rt_sw), 
        .S(top_code_0_n_s_ctrl), .Y(rt_sw_5));
    MX2C dumponoff_rst_RNO_0 (.A(net_33_0), .B(top_code_0_noise_rst_0), 
        .S(top_code_0_n_s_ctrl_0), .Y(dumponoff_rst_5));
    GND GND_i_0 (.Y(GND_0));
    DFN1 dumpon_ctr (.D(dumpon_ctr_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_dumpon_ctr));
    MX2C soft_d_RNO_0 (.A(scanstate_0_soft_d), .B(noisestate_0_soft_d), 
        .S(top_code_0_n_s_ctrl_1), .Y(soft_d_5));
    DFN1 intertodsp (.D(intertodsp_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_intertodsp));
    MX2C dumpon_ctr_RNO_0 (.A(scanstate_0_dds_conf), .B(
        noisestate_0_dumpon_ctr), .S(top_code_0_n_s_ctrl_1), .Y(
        dumpon_ctr_5));
    VCC VCC_i (.Y(VCC));
    NOR2A soft_d_RNO (.A(net_27), .B(soft_d_5), .Y(soft_d_RNO_net_1));
    NOR2A dumpoff_ctr_RNO (.A(net_27), .B(dumpoff_ctr_5), .Y(
        dumpoff_ctr_RNO_net_1));
    NOR2A intertodsp_RNO (.A(net_27), .B(intertodsp_5), .Y(
        intertodsp_RNO_net_1));
    GND GND_i (.Y(GND));
    NOR2A dumponoff_rst_RNO (.A(net_27), .B(dumponoff_rst_5), .Y(
        dumponoff_rst_RNO_net_1));
    OR2B sw_acq2_RNO (.A(sw_acq2_5), .B(net_27), .Y(sw_acq2_RNO_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2A rt_sw_RNO (.A(net_27), .B(rt_sw_5), .Y(rt_sw_RNO_net_1));
    DFN1 dumpoff_ctr (.D(dumpoff_ctr_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_dumpoff_ctr));
    MX2C intertodsp_RNO_0 (.A(scanstate_0_state_over_n), .B(
        noisestate_0_state_over_n), .S(top_code_0_n_s_ctrl_0), .Y(
        intertodsp_5));
    MX2C dumpoff_ctr_RNO_0 (.A(scanstate_0_dumpoff_ctr), .B(
        noisestate_0_dumpoff_ctr), .S(top_code_0_n_s_ctrl_0), .Y(
        dumpoff_ctr_5));
    DFN1 sw_acq2 (.D(sw_acq2_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_sw_acq2));
    DFN1 soft_d (.D(soft_d_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_soft_d));
    DFN1 dumponoff_rst (.D(dumponoff_rst_RNO_net_1), .CLK(GLA), .Q(
        nsctrl_choice_0_dumponoff_rst));
    
endmodule


module scanstate(
       timecount_1_0,
       scandata,
       GLA,
       top_code_0_scanchoice,
       top_code_0_scanload,
       scanstate_0_calctrl,
       scanstate_0_soft_d,
       scanstate_0_dds_conf,
       net_33,
       scanstate_0_state_over_n,
       scanstate_0_s_acq,
       scanstate_0_dumpoff_ctr,
       scanstate_0_rt_sw,
       scanstate_0_sw_acq2,
       net_33_0,
       timer_top_0_clk_en_scan
    );
output [15:0] timecount_1_0;
input  [15:0] scandata;
input  GLA;
input  top_code_0_scanchoice;
input  top_code_0_scanload;
output scanstate_0_calctrl;
output scanstate_0_soft_d;
output scanstate_0_dds_conf;
input  net_33;
output scanstate_0_state_over_n;
output scanstate_0_s_acq;
output scanstate_0_dumpoff_ctr;
output scanstate_0_rt_sw;
output scanstate_0_sw_acq2;
input  net_33_0;
input  timer_top_0_clk_en_scan;

    wire \CS_srsts_i_0[6] , \CS[6]_net_1 , \CS_srsts_i_0[2] , 
        \CS[2]_net_1 , \CS_srsts_i_0[3] , \CS[3]_net_1 , 
        \CS_srsts_i_0[4] , \CS[4]_net_1 , \CS_srsts_i_0[5] , 
        \CS[5]_net_1 , \CS_srsts_i_0[1] , \CS[1]_net_1 , \CS_li[0] , 
        \CS_RNO_0[5]_net_1 , \CS_RNO_0[4]_net_1 , \CS_RNO_0[3]_net_1 , 
        \CS_RNO_0[2]_net_1 , \CS_RNO_0[1]_net_1 , \timecount_cnst[4] , 
        \CS_RNO_0[6]_net_1 , N_114, N_299, N_313, N_116, N_118, N_315, 
        N_63, \acqtime[0]_net_1 , \dectime[0]_net_1 , N_255, N_65, 
        \acqtime[2]_net_1 , \dectime[2]_net_1 , N_67, 
        \acqtime[4]_net_1 , \dectime[4]_net_1 , N_68, 
        \acqtime[5]_net_1 , \dectime[5]_net_1 , N_70, 
        \acqtime[7]_net_1 , \dectime[7]_net_1 , N_71, 
        \acqtime[8]_net_1 , \dectime[8]_net_1 , N_73, 
        \acqtime[10]_net_1 , \dectime[10]_net_1 , N_75, 
        \acqtime[12]_net_1 , \dectime[12]_net_1 , N_76, 
        \acqtime[13]_net_1 , \dectime[13]_net_1 , N_77, 
        \acqtime[14]_net_1 , \dectime[14]_net_1 , N_78, 
        \acqtime[15]_net_1 , \dectime[15]_net_1 , \timecount_5[0] , 
        N_292, \timecount_5[2] , \timecount_cnst[2] , \timecount_5[4] , 
        \timecount_5[5] , \timecount_5[7] , \timecount_5[8] , 
        \timecount_5[10] , \timecount_5[12] , \timecount_5[13] , 
        \timecount_5[14] , \timecount_5[15] , s_acq_RNO_net_1, 
        dumpoff_ctr_RNO_1, rt_sw_RNO_0_net_1, state_over_n_RNO_0, 
        sw_acq2_RNO_0_net_1, \CS_RNO_0[7] , \CS[7]_net_1 , 
        un1_dumpoff_ctr_2_sqmuxa, soft_d_RNO_0_net_1, N_115, 
        dds_conf_RNO_0_net_1, N_136, \CS_i_0_RNO[0]_net_1 , N_249, 
        \timecount_5[11] , N_74, \timecount_5[9] , N_72, 
        \timecount_5[3] , N_66, \acqtime[11]_net_1 , 
        \dectime[11]_net_1 , \acqtime[9]_net_1 , \dectime[9]_net_1 , 
        \acqtime[3]_net_1 , \dectime[3]_net_1 , calctrl_RNO_net_1, 
        N_137, \timecount_5[1] , N_64, \acqtime[1]_net_1 , 
        \dectime[1]_net_1 , \timecount_5[6] , N_69, \acqtime[6]_net_1 , 
        \dectime[6]_net_1 , acqtime_1_sqmuxa_net_1, 
        acqtime_0_sqmuxa_net_1, GND, VCC, GND_0, VCC_0;
    
    DFN1E1 \acqtime[7]  (.D(scandata[7]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[7]_net_1 ));
    MX2C \timecount_1_RNO_0[3]  (.A(\acqtime[3]_net_1 ), .B(
        \dectime[3]_net_1 ), .S(N_255), .Y(N_66));
    MX2C \timecount_1_RNO_0[12]  (.A(\acqtime[12]_net_1 ), .B(
        \dectime[12]_net_1 ), .S(N_255), .Y(N_75));
    NOR2 \timecount_1_RNO[10]  (.A(N_292), .B(N_73), .Y(
        \timecount_5[10] ));
    DFN1E1 \timecount_1[0]  (.D(\timecount_5[0] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[0]));
    DFN1E1 \timecount_1[1]  (.D(\timecount_5[1] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[1]));
    DFN1E1 \dectime[1]  (.D(scandata[1]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[1]_net_1 ));
    DFN1E1 \dectime[2]  (.D(scandata[2]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[2]_net_1 ));
    AO1A calctrl_RNO_0 (.A(\CS[5]_net_1 ), .B(scanstate_0_calctrl), .C(
        \CS[2]_net_1 ), .Y(N_137));
    OA1C \CS_RNO[4]  (.A(timer_top_0_clk_en_scan), .B(\CS[3]_net_1 ), 
        .C(\CS_srsts_i_0[4] ), .Y(\CS_RNO_0[4]_net_1 ));
    OR2A sw_acq2_RNO (.A(net_33), .B(N_114), .Y(sw_acq2_RNO_0_net_1));
    MX2A \timecount_1_RNO[5]  (.A(N_68), .B(net_33_0), .S(N_292), .Y(
        \timecount_5[5] ));
    NOR2B rt_sw_RNO (.A(N_116), .B(net_33_0), .Y(rt_sw_RNO_0_net_1));
    DFN1E1 \acqtime[11]  (.D(scandata[11]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[11]_net_1 ));
    MX2C \timecount_1_RNO[7]  (.A(N_70), .B(\timecount_cnst[4] ), .S(
        N_292), .Y(\timecount_5[7] ));
    OA1 s_acq_RNO (.A(\CS[4]_net_1 ), .B(scanstate_0_s_acq), .C(
        net_33_0), .Y(s_acq_RNO_net_1));
    DFN1 sw_acq2 (.D(sw_acq2_RNO_0_net_1), .CLK(GLA), .Q(
        scanstate_0_sw_acq2));
    DFN1 calctrl (.D(calctrl_RNO_net_1), .CLK(GLA), .Q(
        scanstate_0_calctrl));
    DFN1E1 \acqtime[6]  (.D(scandata[6]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[6]_net_1 ));
    DFN1 \CS[4]  (.D(\CS_RNO_0[4]_net_1 ), .CLK(GLA), .Q(\CS[4]_net_1 )
        );
    DFN1E1 \acqtime[4]  (.D(scandata[4]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[4]_net_1 ));
    DFN1E1 \acqtime[15]  (.D(scandata[15]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[15]_net_1 ));
    OAI1 \CS_RNO_0[4]  (.A(\CS[4]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(net_33_0), .Y(\CS_srsts_i_0[4] ));
    DFN1E1 \timecount_1[13]  (.D(\timecount_5[13] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[13]));
    DFN1E1 \timecount_1[10]  (.D(\timecount_5[10] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[10]));
    MX2C \timecount_1_RNO[6]  (.A(N_69), .B(\timecount_cnst[2] ), .S(
        N_292), .Y(\timecount_5[6] ));
    DFN1E1 \dectime[13]  (.D(scandata[13]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[13]_net_1 ));
    NOR2B acqtime_0_sqmuxa (.A(top_code_0_scanload), .B(
        top_code_0_scanchoice), .Y(acqtime_0_sqmuxa_net_1));
    MX2C \timecount_1_RNO_0[9]  (.A(\acqtime[9]_net_1 ), .B(
        \dectime[9]_net_1 ), .S(N_255), .Y(N_72));
    AO1A dds_conf_RNO_0 (.A(\CS[2]_net_1 ), .B(scanstate_0_dds_conf), 
        .C(\CS[1]_net_1 ), .Y(N_136));
    DFN1E1 \dectime[10]  (.D(scandata[10]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[10]_net_1 ));
    DFN1E1 \timecount_1[2]  (.D(\timecount_5[2] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[2]));
    MX2 soft_d_RNO_0 (.A(scanstate_0_soft_d), .B(\CS[1]_net_1 ), .S(
        N_313), .Y(N_115));
    DFN1 \CS_i_0[0]  (.D(\CS_i_0_RNO[0]_net_1 ), .CLK(GLA), .Q(
        \CS_li[0] ));
    DFN1 \CS[3]  (.D(\CS_RNO_0[3]_net_1 ), .CLK(GLA), .Q(\CS[3]_net_1 )
        );
    OR2B \CS_RNI1AU9[1]  (.A(\CS[1]_net_1 ), .B(net_33), .Y(N_249));
    DFN1E1 \timecount_1[12]  (.D(\timecount_5[12] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[12]));
    DFN1E1 \dectime[8]  (.D(scandata[8]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[8]_net_1 ));
    OA1C \CS_RNO[5]  (.A(timer_top_0_clk_en_scan), .B(\CS[4]_net_1 ), 
        .C(\CS_srsts_i_0[5] ), .Y(\CS_RNO_0[5]_net_1 ));
    OAI1 \CS_RNO_0[5]  (.A(\CS[5]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(net_33_0), .Y(\CS_srsts_i_0[5] ));
    MX2C \timecount_1_RNO_0[5]  (.A(\acqtime[5]_net_1 ), .B(
        \dectime[5]_net_1 ), .S(N_255), .Y(N_68));
    NOR2B dumpoff_ctr_RNO (.A(N_118), .B(net_33_0), .Y(
        dumpoff_ctr_RNO_1));
    MX2A \CS_RNO_0[1]  (.A(\CS[1]_net_1 ), .B(\CS_li[0] ), .S(
        timer_top_0_clk_en_scan), .Y(\CS_srsts_i_0[1] ));
    DFN1E1 \acqtime[10]  (.D(scandata[10]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[10]_net_1 ));
    DFN1E1 \timecount_1[8]  (.D(\timecount_5[8] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[8]));
    MX2C \timecount_1_RNO_0[10]  (.A(\acqtime[10]_net_1 ), .B(
        \dectime[10]_net_1 ), .S(N_255), .Y(N_73));
    DFN1 \CS[1]  (.D(\CS_RNO_0[1]_net_1 ), .CLK(GLA), .Q(\CS[1]_net_1 )
        );
    GND GND_i (.Y(GND));
    DFN1E1 \dectime[15]  (.D(scandata[15]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[15]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    MX2C \timecount_1_RNO_0[4]  (.A(\acqtime[4]_net_1 ), .B(
        \dectime[4]_net_1 ), .S(N_255), .Y(N_67));
    MX2C \timecount_1_RNO_0[2]  (.A(\acqtime[2]_net_1 ), .B(
        \dectime[2]_net_1 ), .S(N_255), .Y(N_65));
    OA1B \CS_RNO[7]  (.A(\CS[7]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(un1_dumpoff_ctr_2_sqmuxa), .Y(\CS_RNO_0[7] ));
    MX2C \timecount_1_RNO[4]  (.A(N_67), .B(\timecount_cnst[4] ), .S(
        N_292), .Y(\timecount_5[4] ));
    DFN1E1 \timecount_1[11]  (.D(\timecount_5[11] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[11]));
    NOR2B soft_d_RNO (.A(N_115), .B(net_33), .Y(soft_d_RNO_0_net_1));
    DFN1E1 \acqtime[14]  (.D(scandata[14]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[14]_net_1 ));
    DFN1E1 \timecount_1[5]  (.D(\timecount_5[5] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[5]));
    OA1C \CS_RNO[3]  (.A(timer_top_0_clk_en_scan), .B(\CS[2]_net_1 ), 
        .C(\CS_srsts_i_0[3] ), .Y(\CS_RNO_0[3]_net_1 ));
    DFN1E1 \timecount_1[14]  (.D(\timecount_5[14] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[14]));
    DFN1 soft_d (.D(soft_d_RNO_0_net_1), .CLK(GLA), .Q(
        scanstate_0_soft_d));
    DFN1E1 \acqtime[9]  (.D(scandata[9]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[9]_net_1 ));
    NOR2 \CS_RNIJQBB[6]  (.A(\CS[7]_net_1 ), .B(\CS[6]_net_1 ), .Y(
        N_315));
    OAI1 \CS_RNO_0[6]  (.A(\CS[6]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(net_33_0), .Y(\CS_srsts_i_0[6] ));
    OA1 \CS_i_0_RNO[0]  (.A(\CS_li[0] ), .B(timer_top_0_clk_en_scan), 
        .C(net_33), .Y(\CS_i_0_RNO[0]_net_1 ));
    DFN1 state_over_n (.D(state_over_n_RNO_0), .CLK(GLA), .Q(
        scanstate_0_state_over_n));
    NOR2A \CS_RNO[1]  (.A(net_33_0), .B(\CS_srsts_i_0[1] ), .Y(
        \CS_RNO_0[1]_net_1 ));
    MX2C \timecount_1_RNO[3]  (.A(N_66), .B(N_249), .S(N_292), .Y(
        \timecount_5[3] ));
    NOR2B dds_conf_RNO (.A(N_136), .B(net_33), .Y(dds_conf_RNO_0_net_1)
        );
    VCC VCC_i (.Y(VCC));
    DFN1E1 \timecount_1[7]  (.D(\timecount_5[7] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[7]));
    DFN1E1 \dectime[12]  (.D(scandata[12]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[12]_net_1 ));
    OAI1 \CS_RNO_0[2]  (.A(\CS[2]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(net_33_0), .Y(\CS_srsts_i_0[2] ));
    DFN1E1 \acqtime[2]  (.D(scandata[2]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[2]_net_1 ));
    NOR2 \timecount_1_RNO[12]  (.A(N_292), .B(N_75), .Y(
        \timecount_5[12] ));
    MX2B rt_sw_RNO_0 (.A(scanstate_0_rt_sw), .B(\CS[5]_net_1 ), .S(
        N_313), .Y(N_116));
    OR3B \CS_i_0_RNI3J7C[0]  (.A(\CS_li[0] ), .B(net_33_0), .C(
        \CS[5]_net_1 ), .Y(\timecount_cnst[4] ));
    DFN1E1 \timecount_1[15]  (.D(\timecount_5[15] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[15]));
    OAI1 \CS_RNIFCEH[2]  (.A(\CS[2]_net_1 ), .B(\CS[4]_net_1 ), .C(
        net_33_0), .Y(N_292));
    DFN1E1 \dectime[6]  (.D(scandata[6]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[6]_net_1 ));
    DFN1 dumpoff_ctr (.D(dumpoff_ctr_RNO_1), .CLK(GLA), .Q(
        scanstate_0_dumpoff_ctr));
    MX2C \timecount_1_RNO_0[1]  (.A(\acqtime[1]_net_1 ), .B(
        \dectime[1]_net_1 ), .S(N_255), .Y(N_64));
    NOR2B \CS_i_0_RNIBUQB[0]  (.A(N_315), .B(\CS_li[0] ), .Y(N_313));
    MX2C \timecount_1_RNO_0[13]  (.A(\acqtime[13]_net_1 ), .B(
        \dectime[13]_net_1 ), .S(N_255), .Y(N_76));
    MX2C \timecount_1_RNO_0[11]  (.A(\acqtime[11]_net_1 ), .B(
        \dectime[11]_net_1 ), .S(N_255), .Y(N_74));
    MX2C \timecount_1_RNO[0]  (.A(N_63), .B(net_33_0), .S(N_292), .Y(
        \timecount_5[0] ));
    DFN1E1 \timecount_1[6]  (.D(\timecount_5[6] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[6]));
    NOR2 sw_acq2_RNO_1 (.A(\CS[4]_net_1 ), .B(\CS[3]_net_1 ), .Y(N_299)
        );
    DFN1 \CS[7]  (.D(\CS_RNO_0[7] ), .CLK(GLA), .Q(\CS[7]_net_1 ));
    NOR2 \timecount_1_RNO[15]  (.A(N_292), .B(N_78), .Y(
        \timecount_5[15] ));
    DFN1 s_acq (.D(s_acq_RNO_net_1), .CLK(GLA), .Q(scanstate_0_s_acq));
    DFN1 \CS[6]  (.D(\CS_RNO_0[6]_net_1 ), .CLK(GLA), .Q(\CS[6]_net_1 )
        );
    DFN1E1 \dectime[0]  (.D(scandata[0]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[0]_net_1 ));
    AO1B state_over_n_RNO (.A(scanstate_0_state_over_n), .B(N_315), .C(
        net_33), .Y(state_over_n_RNO_0));
    MX2C \timecount_1_RNO_0[0]  (.A(\acqtime[0]_net_1 ), .B(
        \dectime[0]_net_1 ), .S(N_255), .Y(N_63));
    DFN1E1 \acqtime[1]  (.D(scandata[1]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[1]_net_1 ));
    MX2C \timecount_1_RNO_0[6]  (.A(\acqtime[6]_net_1 ), .B(
        \dectime[6]_net_1 ), .S(N_255), .Y(N_69));
    OA1C \CS_RNO[2]  (.A(timer_top_0_clk_en_scan), .B(\CS[1]_net_1 ), 
        .C(\CS_srsts_i_0[2] ), .Y(\CS_RNO_0[2]_net_1 ));
    GND GND_i_0 (.Y(GND_0));
    MX2C \timecount_1_RNO_0[8]  (.A(\acqtime[8]_net_1 ), .B(
        \dectime[8]_net_1 ), .S(N_255), .Y(N_71));
    DFN1E1 \acqtime[0]  (.D(scandata[0]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[0]_net_1 ));
    NOR2 \timecount_1_RNO[1]  (.A(N_292), .B(N_64), .Y(
        \timecount_5[1] ));
    OR2A \CS_RNI1AU9_0[1]  (.A(net_33), .B(\CS[1]_net_1 ), .Y(
        \timecount_cnst[2] ));
    MX2 sw_acq2_RNO_0 (.A(scanstate_0_sw_acq2), .B(N_299), .S(N_313), 
        .Y(N_114));
    AO1 dumpoff_ctr_RNO_0 (.A(scanstate_0_dumpoff_ctr), .B(N_315), .C(
        \CS[5]_net_1 ), .Y(N_118));
    DFN1E1 \acqtime[8]  (.D(scandata[8]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[8]_net_1 ));
    OR2A \CS_RNIG7KF[6]  (.A(net_33), .B(N_315), .Y(
        un1_dumpoff_ctr_2_sqmuxa));
    DFN1 \CS[2]  (.D(\CS_RNO_0[2]_net_1 ), .CLK(GLA), .Q(\CS[2]_net_1 )
        );
    DFN1E1 \dectime[11]  (.D(scandata[11]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[11]_net_1 ));
    DFN1E1 \dectime[4]  (.D(scandata[4]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[4]_net_1 ));
    NOR2 \timecount_1_RNO[13]  (.A(N_292), .B(N_76), .Y(
        \timecount_5[13] ));
    DFN1E1 \acqtime[5]  (.D(scandata[5]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[5]_net_1 ));
    DFN1 dds_conf (.D(dds_conf_RNO_0_net_1), .CLK(GLA), .Q(
        scanstate_0_dds_conf));
    DFN1E1 \timecount_1[9]  (.D(\timecount_5[9] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[9]));
    DFN1E1 \dectime[3]  (.D(scandata[3]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[3]_net_1 ));
    NOR2 \timecount_1_RNO[14]  (.A(N_292), .B(N_77), .Y(
        \timecount_5[14] ));
    DFN1 \CS[5]  (.D(\CS_RNO_0[5]_net_1 ), .CLK(GLA), .Q(\CS[5]_net_1 )
        );
    MX2C \timecount_1_RNO[2]  (.A(N_65), .B(\timecount_cnst[2] ), .S(
        N_292), .Y(\timecount_5[2] ));
    OAI1 \CS_RNO_0[3]  (.A(\CS[3]_net_1 ), .B(timer_top_0_clk_en_scan), 
        .C(net_33_0), .Y(\CS_srsts_i_0[3] ));
    DFN1E1 \acqtime[3]  (.D(scandata[3]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[3]_net_1 ));
    DFN1E1 \timecount_1[3]  (.D(\timecount_5[3] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[3]));
    MX2C \timecount_1_RNO[9]  (.A(N_72), .B(N_249), .S(N_292), .Y(
        \timecount_5[9] ));
    DFN1 rt_sw (.D(rt_sw_RNO_0_net_1), .CLK(GLA), .Q(scanstate_0_rt_sw)
        );
    DFN1E1 \dectime[14]  (.D(scandata[14]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[14]_net_1 ));
    DFN1E1 \dectime[7]  (.D(scandata[7]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[7]_net_1 ));
    OA1C \CS_RNO[6]  (.A(timer_top_0_clk_en_scan), .B(\CS[5]_net_1 ), 
        .C(\CS_srsts_i_0[6] ), .Y(\CS_RNO_0[6]_net_1 ));
    NOR2B calctrl_RNO (.A(N_137), .B(net_33), .Y(calctrl_RNO_net_1));
    MX2C \timecount_1_RNO[11]  (.A(N_74), .B(N_249), .S(N_292), .Y(
        \timecount_5[11] ));
    MX2C \timecount_1_RNO_0[7]  (.A(\acqtime[7]_net_1 ), .B(
        \dectime[7]_net_1 ), .S(N_255), .Y(N_70));
    OR2B \CS_RNI4AU9[4]  (.A(\CS[4]_net_1 ), .B(net_33), .Y(N_255));
    MX2C \timecount_1_RNO[8]  (.A(N_71), .B(\timecount_cnst[4] ), .S(
        N_292), .Y(\timecount_5[8] ));
    DFN1E1 \dectime[9]  (.D(scandata[9]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[9]_net_1 ));
    DFN1E1 \acqtime[13]  (.D(scandata[13]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[13]_net_1 ));
    DFN1E1 \acqtime[12]  (.D(scandata[12]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[12]_net_1 ));
    DFN1E1 \timecount_1[4]  (.D(\timecount_5[4] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1_0[4]));
    DFN1E1 \dectime[5]  (.D(scandata[5]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[5]_net_1 ));
    MX2C \timecount_1_RNO_0[15]  (.A(\acqtime[15]_net_1 ), .B(
        \dectime[15]_net_1 ), .S(N_255), .Y(N_78));
    NOR2A acqtime_1_sqmuxa (.A(top_code_0_scanload), .B(
        top_code_0_scanchoice), .Y(acqtime_1_sqmuxa_net_1));
    MX2C \timecount_1_RNO_0[14]  (.A(\acqtime[14]_net_1 ), .B(
        \dectime[14]_net_1 ), .S(N_255), .Y(N_77));
    
endmodule


module off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1(
       i_3,
       GLA,
       DUMP_OFF_0_dump_off,
       off_on_state_0_state_over,
       bri_dump_sw_0_reset_out_0
    );
input  [1:0] i_3;
input  GLA;
output DUMP_OFF_0_dump_off;
output off_on_state_0_state_over;
input  bri_dump_sw_0_reset_out_0;

    wire N_14, N_13, N_42, \cs_ns[1] , \cs[1]_net_1 , \cs_nsss[1] , 
        \cs_nsss[0] , GND, VCC, GND_0, VCC_0;
    
    OR2B state_over_RNO_0 (.A(off_on_state_0_state_over), .B(N_42), .Y(
        N_13));
    DFN1 state_over (.D(N_14), .CLK(GLA), .Q(off_on_state_0_state_over)
        );
    DFN1 \cs[0]  (.D(\cs_nsss[0] ), .CLK(GLA), .Q(DUMP_OFF_0_dump_off));
    NOR3C \cs_RNO[0]  (.A(N_42), .B(bri_dump_sw_0_reset_out_0), .C(
        i_3[0]), .Y(\cs_nsss[0] ));
    VCC VCC_i_0 (.Y(VCC_0));
    DFN1 \cs[1]  (.D(\cs_nsss[1] ), .CLK(GLA), .Q(\cs[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3C \cs_RNO[1]  (.A(\cs_ns[1] ), .B(bri_dump_sw_0_reset_out_0), 
        .C(i_3[0]), .Y(\cs_nsss[1] ));
    AOI1 \cs_RNIIT8E[1]  (.A(DUMP_OFF_0_dump_off), .B(i_3[1]), .C(
        \cs[1]_net_1 ), .Y(N_42));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    MX2 \cs_RNO_0[1]  (.A(\cs[1]_net_1 ), .B(i_3[1]), .S(
        DUMP_OFF_0_dump_off), .Y(\cs_ns[1] ));
    OR3C state_over_RNO (.A(N_13), .B(i_3[0]), .C(
        bri_dump_sw_0_reset_out_0), .Y(N_14));
    
endmodule


module off_on_coder(
       i_3,
       count_3,
       GLA,
       bri_dump_sw_0_dumpoff_ctr,
       bri_dump_sw_0_reset_out_0
    );
output [1:0] i_3;
input  [4:0] count_3;
input  GLA;
input  bri_dump_sw_0_dumpoff_ctr;
input  bri_dump_sw_0_reset_out_0;

    wire \i_0_1[1] , \i_RNO_1[1]_net_1 , N_17, \i_RNO_0[0] , GND, VCC, 
        GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2 \i_RNO_1[1]  (.A(count_3[1]), .B(count_3[0]), .Y(N_17));
    DFN1 \i[1]  (.D(\i_RNO_1[1]_net_1 ), .CLK(GLA), .Q(i_3[1]));
    GND GND_i_0 (.Y(GND_0));
    NOR3C \i_RNO[1]  (.A(\i_0_1[1] ), .B(N_17), .C(
        bri_dump_sw_0_reset_out_0), .Y(\i_RNO_1[1]_net_1 ));
    VCC VCC_i (.Y(VCC));
    NOR3B \i_RNO_0[1]  (.A(count_3[2]), .B(count_3[4]), .C(count_3[3]), 
        .Y(\i_0_1[1] ));
    NOR2B \i_RNO[0]  (.A(bri_dump_sw_0_reset_out_0), .B(
        bri_dump_sw_0_dumpoff_ctr), .Y(\i_RNO_0[0] ));
    DFN1 \i[0]  (.D(\i_RNO_0[0] ), .CLK(GLA), .Q(i_3[0]));
    GND GND_i (.Y(GND));
    
endmodule


module off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0(
       count_3,
       GLA,
       bri_dump_sw_0_reset_out_0,
       off_on_state_0_state_over,
       bri_dump_sw_0_dumpoff_ctr
    );
output [4:0] count_3;
input  GLA;
input  bri_dump_sw_0_reset_out_0;
input  off_on_state_0_state_over;
input  bri_dump_sw_0_dumpoff_ctr;

    wire N_5, count_0_sqmuxa_net_1, N_7, N_12, N_9, N_13, count_n0, 
        N_11, N_14, GND, VCC, GND_0, VCC_0;
    
    NOR2B \count_RNI9785[1]  (.A(count_3[1]), .B(count_3[0]), .Y(N_12));
    GND GND_i_0 (.Y(GND_0));
    XA1B \count_RNO[1]  (.A(count_3[0]), .B(count_3[1]), .C(
        count_0_sqmuxa_net_1), .Y(N_5));
    DFN1 \count[3]  (.D(N_9), .CLK(GLA), .Q(count_3[3]));
    DFN1 \count[0]  (.D(count_n0), .CLK(GLA), .Q(count_3[0]));
    XA1B \count_RNO[3]  (.A(N_13), .B(count_3[3]), .C(
        count_0_sqmuxa_net_1), .Y(N_9));
    NOR2B \count_RNIVGS7[2]  (.A(count_3[2]), .B(N_12), .Y(N_13));
    VCC VCC_i (.Y(VCC));
    GND GND_i (.Y(GND));
    NOR2B \count_RNO_0[4]  (.A(count_3[3]), .B(N_13), .Y(N_14));
    XA1B \count_RNO[2]  (.A(N_12), .B(count_3[2]), .C(
        count_0_sqmuxa_net_1), .Y(N_7));
    OR3C count_0_sqmuxa (.A(bri_dump_sw_0_dumpoff_ctr), .B(
        off_on_state_0_state_over), .C(bri_dump_sw_0_reset_out_0), .Y(
        count_0_sqmuxa_net_1));
    VCC VCC_i_0 (.Y(VCC_0));
    XA1B \count_RNO[4]  (.A(N_14), .B(count_3[4]), .C(
        count_0_sqmuxa_net_1), .Y(N_11));
    DFN1 \count[1]  (.D(N_5), .CLK(GLA), .Q(count_3[1]));
    DFN1 \count[4]  (.D(N_11), .CLK(GLA), .Q(count_3[4]));
    NOR2 \count_RNO[0]  (.A(count_3[0]), .B(count_0_sqmuxa_net_1), .Y(
        count_n0));
    DFN1 \count[2]  (.D(N_7), .CLK(GLA), .Q(count_3[2]));
    
endmodule


module DUMP_OFF_DUMP_OFF_0(
       bri_dump_sw_0_dumpoff_ctr,
       bri_dump_sw_0_reset_out_0,
       DUMP_OFF_0_dump_off,
       GLA
    );
input  bri_dump_sw_0_dumpoff_ctr;
input  bri_dump_sw_0_reset_out_0;
output DUMP_OFF_0_dump_off;
input  GLA;

    wire \i_3[0] , \i_3[1] , off_on_state_0_state_over, \count_3[0] , 
        \count_3[1] , \count_3[2] , \count_3[3] , \count_3[4] , GND, 
        VCC, GND_0, VCC_0;
    
    VCC VCC_i_0 (.Y(VCC_0));
    off_on_state_DUMP_0_off_on_state_1_DUMP_0_off_on_state_1 
        off_on_state_0 (.i_3({\i_3[1] , \i_3[0] }), .GLA(GLA), 
        .DUMP_OFF_0_dump_off(DUMP_OFF_0_dump_off), 
        .off_on_state_0_state_over(off_on_state_0_state_over), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0));
    off_on_coder off_on_coder_0 (.i_3({\i_3[1] , \i_3[0] }), .count_3({
        \count_3[4] , \count_3[3] , \count_3[2] , \count_3[1] , 
        \count_3[0] }), .GLA(GLA), .bri_dump_sw_0_dumpoff_ctr(
        bri_dump_sw_0_dumpoff_ctr), .bri_dump_sw_0_reset_out_0(
        bri_dump_sw_0_reset_out_0));
    GND GND_i_0 (.Y(GND_0));
    VCC VCC_i (.Y(VCC));
    off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0 
        off_on_timer_0 (.count_3({\count_3[4] , \count_3[3] , 
        \count_3[2] , \count_3[1] , \count_3[0] }), .GLA(GLA), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), 
        .off_on_state_0_state_over(off_on_state_0_state_over), 
        .bri_dump_sw_0_dumpoff_ctr(bri_dump_sw_0_dumpoff_ctr));
    GND GND_i (.Y(GND));
    
endmodule


module n_pluse_acq(
       n_acq_change_0_n_acq_start,
       n_acq_change_0_n_rst_n,
       net_27,
       noisestate_0_n_acq,
       plusestate_0_pluse_acq,
       top_code_0_pluse_noise_ctrl,
       top_code_0_noise_rst_0,
       top_code_0_pluse_rst,
       GLA,
       n_acq_change_0_n_rst_n_0
    );
output n_acq_change_0_n_acq_start;
output n_acq_change_0_n_rst_n;
input  net_27;
input  noisestate_0_n_acq;
input  plusestate_0_pluse_acq;
input  top_code_0_pluse_noise_ctrl;
input  top_code_0_noise_rst_0;
input  top_code_0_pluse_rst;
input  GLA;
output n_acq_change_0_n_rst_n_0;

    wire n_rst_n_0_net_1, n_rst_n_5_net_1, n_acq_start_5, 
        n_acq_start_RNO_net_1, GND, VCC, GND_0, VCC_0;
    
    NOR2A n_rst_n_0 (.A(net_27), .B(n_rst_n_5_net_1), .Y(
        n_rst_n_0_net_1));
    DFN1 n_acq_start (.D(n_acq_start_RNO_net_1), .CLK(GLA), .Q(
        n_acq_change_0_n_acq_start));
    MX2C n_rst_n_5 (.A(top_code_0_pluse_rst), .B(
        top_code_0_noise_rst_0), .S(top_code_0_pluse_noise_ctrl), .Y(
        n_rst_n_5_net_1));
    DFN1 n_rst_n (.D(n_rst_n_0_net_1), .CLK(GLA), .Q(
        n_acq_change_0_n_rst_n));
    VCC VCC_i_0 (.Y(VCC_0));
    NOR2A n_acq_start_RNO (.A(net_27), .B(n_acq_start_5), .Y(
        n_acq_start_RNO_net_1));
    VCC VCC_i (.Y(VCC));
    DFN1 n_rst_n_0_0 (.D(n_rst_n_0_net_1), .CLK(GLA), .Q(
        n_acq_change_0_n_rst_n_0));
    MX2C n_acq_start_RNO_0 (.A(plusestate_0_pluse_acq), .B(
        noisestate_0_n_acq), .S(top_code_0_pluse_noise_ctrl), .Y(
        n_acq_start_5));
    GND GND_i_0 (.Y(GND_0));
    GND GND_i (.Y(GND));
    
endmodule


module noisestate(
       timecount_1,
       noisedata,
       GLA,
       noisestate_0_soft_d,
       noisestate_0_sw_acq2,
       noisestate_0_rt_sw,
       noisestate_0_n_acq,
       top_code_0_nstatechoice,
       top_code_0_nstateload,
       noisestate_0_dumpoff_ctr,
       top_code_0_noise_rst,
       noisestate_0_dumpon_ctr,
       noisestate_0_state_over_n,
       top_code_0_noise_rst_0,
       timer_top_0_clk_en_noise
    );
output [15:0] timecount_1;
input  [15:0] noisedata;
input  GLA;
output noisestate_0_soft_d;
output noisestate_0_sw_acq2;
output noisestate_0_rt_sw;
output noisestate_0_n_acq;
input  top_code_0_nstatechoice;
input  top_code_0_nstateload;
output noisestate_0_dumpoff_ctr;
input  top_code_0_noise_rst;
output noisestate_0_dumpon_ctr;
output noisestate_0_state_over_n;
input  top_code_0_noise_rst_0;
input  timer_top_0_clk_en_noise;

    wire \CS_srsts_i_0[2] , \CS[2]_net_1 , \CS_srsts_i_0[3] , 
        \CS[3]_net_1 , \CS_srsts_i_0[4] , \CS[4]_net_1 , 
        \CS_srsts_i_0[6] , \CS[6]_net_1 , \CS_srsts_i_0[1] , 
        \CS[1]_net_1 , \CS_li[0] , \CS_RNO_2[6] , \CS[5]_net_1 , 
        \CS_RNO_2[5] , N_296, N_295, \CS_RNO_2[4] , \CS_RNO_2[3] , 
        \timecount_cnst[4] , \CS_RNO_2[1] , \CS_RNO_2[2] , 
        \timecount_5[7] , N_68, N_280, state_over_n_RNO_1, N_302, 
        dumpon_ctr_RNO_0_net_1, N_134, N_282, \timecount_5[11] , N_72, 
        N_243, \timecount_5[9] , N_70, \timecount_5[3] , N_64, 
        \acqtime[11]_net_1 , \dectime[11]_net_1 , N_245, 
        \acqtime[9]_net_1 , \dectime[9]_net_1 , \acqtime[3]_net_1 , 
        \dectime[3]_net_1 , \CS_RNO_2[7] , \CS[7]_net_1 , 
        un1_dumpoff_ctr_2_sqmuxa, dumpoff_ctr_RNO_2, N_116, N_300, 
        \timecount_5[8] , N_69, \timecount_5[4] , N_65, 
        \dectime[8]_net_1 , \acqtime[8]_net_1 , \dectime[4]_net_1 , 
        \acqtime[4]_net_1 , N_63, \dectime[2]_net_1 , 
        \acqtime[2]_net_1 , N_74, \dectime[13]_net_1 , 
        \acqtime[13]_net_1 , \timecount_5[13] , \CS_i_0_RNO_0[0] , 
        acqtime_1_sqmuxa_net_1, acqtime_0_sqmuxa_net_1, 
        sw_acq2_RNO_1_net_1, N_112, rt_sw_RNO_2, N_114, 
        n_acq_RNO_net_1, N_133, N_286, \acqtime[7]_net_1 , 
        \dectime[7]_net_1 , \timecount_5[2] , \timecount_cnst[2] , 
        N_113, soft_d_RNO_1, \timecount_5[15] , N_76, 
        \timecount_5[14] , N_75, \timecount_5[12] , N_73, 
        \timecount_5[10] , N_71, \timecount_5[1] , N_62, 
        \timecount_5[6] , N_67, \timecount_5[5] , N_66, 
        \timecount_5[0] , N_61, \acqtime[15]_net_1 , 
        \dectime[15]_net_1 , \acqtime[14]_net_1 , \dectime[14]_net_1 , 
        \acqtime[12]_net_1 , \dectime[12]_net_1 , \acqtime[10]_net_1 , 
        \dectime[10]_net_1 , \acqtime[6]_net_1 , \dectime[6]_net_1 , 
        \acqtime[5]_net_1 , \dectime[5]_net_1 , \acqtime[1]_net_1 , 
        \dectime[1]_net_1 , \acqtime[0]_net_1 , \dectime[0]_net_1 , 
        GND, VCC, GND_0, VCC_0;
    
    DFN1E1 \acqtime[7]  (.D(noisedata[7]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[7]_net_1 ));
    MX2 \timecount_1_RNO_0[3]  (.A(\acqtime[3]_net_1 ), .B(
        \dectime[3]_net_1 ), .S(N_245), .Y(N_64));
    MX2C \timecount_1_RNO_0[12]  (.A(\acqtime[12]_net_1 ), .B(
        \dectime[12]_net_1 ), .S(N_245), .Y(N_73));
    NOR2 \timecount_1_RNO[10]  (.A(N_280), .B(N_71), .Y(
        \timecount_5[10] ));
    DFN1E1 \timecount_1[0]  (.D(\timecount_5[0] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[0]));
    DFN1E1 \timecount_1[1]  (.D(\timecount_5[1] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[1]));
    DFN1E1 \dectime[1]  (.D(noisedata[1]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[1]_net_1 ));
    DFN1E1 \dectime[2]  (.D(noisedata[2]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[2]_net_1 ));
    OA1C \CS_RNO[4]  (.A(timer_top_0_clk_en_noise), .B(\CS[3]_net_1 ), 
        .C(\CS_srsts_i_0[4] ), .Y(\CS_RNO_2[4] ));
    OR2A sw_acq2_RNO (.A(top_code_0_noise_rst), .B(N_112), .Y(
        sw_acq2_RNO_1_net_1));
    MX2A \timecount_1_RNO[5]  (.A(N_66), .B(top_code_0_noise_rst), .S(
        N_280), .Y(\timecount_5[5] ));
    NOR2B rt_sw_RNO (.A(top_code_0_noise_rst), .B(N_114), .Y(
        rt_sw_RNO_2));
    DFN1E1 \acqtime[11]  (.D(noisedata[11]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[11]_net_1 ));
    MX2C \timecount_1_RNO[7]  (.A(N_68), .B(\timecount_cnst[4] ), .S(
        N_280), .Y(\timecount_5[7] ));
    DFN1 sw_acq2 (.D(sw_acq2_RNO_1_net_1), .CLK(GLA), .Q(
        noisestate_0_sw_acq2));
    DFN1E1 \acqtime[6]  (.D(noisedata[6]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[6]_net_1 ));
    DFN1 \CS[4]  (.D(\CS_RNO_2[4] ), .CLK(GLA), .Q(\CS[4]_net_1 ));
    DFN1E1 \acqtime[4]  (.D(noisedata[4]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[4]_net_1 ));
    DFN1E1 \acqtime[15]  (.D(noisedata[15]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[15]_net_1 ));
    OR2A \CS_RNI1CQA[1]  (.A(top_code_0_noise_rst), .B(\CS[1]_net_1 ), 
        .Y(\timecount_cnst[2] ));
    OAI1 \CS_RNO_0[4]  (.A(\CS[4]_net_1 ), .B(timer_top_0_clk_en_noise)
        , .C(top_code_0_noise_rst_0), .Y(\CS_srsts_i_0[4] ));
    DFN1E1 \timecount_1[13]  (.D(\timecount_5[13] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[13]));
    NOR2B dumpon_ctr_RNO (.A(top_code_0_noise_rst_0), .B(N_134), .Y(
        dumpon_ctr_RNO_0_net_1));
    DFN1E1 \timecount_1[10]  (.D(\timecount_5[10] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[10]));
    MX2C \timecount_1_RNO[6]  (.A(N_67), .B(\timecount_cnst[2] ), .S(
        N_280), .Y(\timecount_5[6] ));
    DFN1E1 \dectime[13]  (.D(noisedata[13]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[13]_net_1 ));
    NOR2B acqtime_0_sqmuxa (.A(top_code_0_nstateload), .B(
        top_code_0_nstatechoice), .Y(acqtime_0_sqmuxa_net_1));
    MX2 \timecount_1_RNO_0[9]  (.A(\acqtime[9]_net_1 ), .B(
        \dectime[9]_net_1 ), .S(N_245), .Y(N_70));
    DFN1E1 \dectime[10]  (.D(noisedata[10]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[10]_net_1 ));
    DFN1E1 \timecount_1[2]  (.D(\timecount_5[2] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[2]));
    MX2 soft_d_RNO_0 (.A(noisestate_0_soft_d), .B(\CS[1]_net_1 ), .S(
        N_300), .Y(N_113));
    DFN1 \CS_i_0[0]  (.D(\CS_i_0_RNO_0[0] ), .CLK(GLA), .Q(\CS_li[0] ));
    DFN1 \CS[3]  (.D(\CS_RNO_2[3] ), .CLK(GLA), .Q(\CS[3]_net_1 ));
    DFN1E1 \timecount_1[12]  (.D(\timecount_5[12] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[12]));
    DFN1E1 \dectime[8]  (.D(noisedata[8]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[8]_net_1 ));
    NOR3A \CS_RNO[5]  (.A(top_code_0_noise_rst_0), .B(N_296), .C(N_295)
        , .Y(\CS_RNO_2[5] ));
    NOR2 \CS_RNO_0[5]  (.A(timer_top_0_clk_en_noise), .B(\CS[5]_net_1 )
        , .Y(N_296));
    MX2C \timecount_1_RNO_0[5]  (.A(\acqtime[5]_net_1 ), .B(
        \dectime[5]_net_1 ), .S(N_245), .Y(N_66));
    NOR2B dumpoff_ctr_RNO (.A(top_code_0_noise_rst_0), .B(N_116), .Y(
        dumpoff_ctr_RNO_2));
    MX2A \CS_RNO_0[1]  (.A(\CS[1]_net_1 ), .B(\CS_li[0] ), .S(
        timer_top_0_clk_en_noise), .Y(\CS_srsts_i_0[1] ));
    DFN1E1 \acqtime[10]  (.D(noisedata[10]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[10]_net_1 ));
    DFN1E1 \timecount_1[8]  (.D(\timecount_5[8] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[8]));
    MX2C \timecount_1_RNO_0[10]  (.A(\acqtime[10]_net_1 ), .B(
        \dectime[10]_net_1 ), .S(N_245), .Y(N_71));
    DFN1 \CS[1]  (.D(\CS_RNO_2[1] ), .CLK(GLA), .Q(\CS[1]_net_1 ));
    GND GND_i (.Y(GND));
    DFN1E1 \dectime[15]  (.D(noisedata[15]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[15]_net_1 ));
    VCC VCC_i_0 (.Y(VCC_0));
    MX2C \timecount_1_RNO_0[4]  (.A(\dectime[4]_net_1 ), .B(
        \acqtime[4]_net_1 ), .S(\CS[4]_net_1 ), .Y(N_65));
    MX2C \timecount_1_RNO_0[2]  (.A(\dectime[2]_net_1 ), .B(
        \acqtime[2]_net_1 ), .S(\CS[4]_net_1 ), .Y(N_63));
    OA1B \CS_RNO[7]  (.A(\CS[7]_net_1 ), .B(timer_top_0_clk_en_noise), 
        .C(un1_dumpoff_ctr_2_sqmuxa), .Y(\CS_RNO_2[7] ));
    MX2C \timecount_1_RNO[4]  (.A(N_65), .B(\timecount_cnst[4] ), .S(
        N_280), .Y(\timecount_5[4] ));
    DFN1E1 \timecount_1[11]  (.D(\timecount_5[11] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[11]));
    NOR2B soft_d_RNO (.A(top_code_0_noise_rst), .B(N_113), .Y(
        soft_d_RNO_1));
    MX2 dumpon_ctr_RNO_0 (.A(N_243), .B(noisestate_0_dumpon_ctr), .S(
        N_282), .Y(N_134));
    DFN1E1 \acqtime[14]  (.D(noisedata[14]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[14]_net_1 ));
    NOR2B \CS_i_0_RNICR9D[0]  (.A(N_302), .B(\CS_li[0] ), .Y(N_300));
    DFN1E1 \timecount_1[5]  (.D(\timecount_5[5] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[5]));
    OA1C \CS_RNO[3]  (.A(timer_top_0_clk_en_noise), .B(\CS[2]_net_1 ), 
        .C(\CS_srsts_i_0[3] ), .Y(\CS_RNO_2[3] ));
    DFN1E1 \timecount_1[14]  (.D(\timecount_5[14] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[14]));
    DFN1 soft_d (.D(soft_d_RNO_1), .CLK(GLA), .Q(noisestate_0_soft_d));
    NOR2 dumpon_ctr_RNO_1 (.A(\CS[2]_net_1 ), .B(\CS[1]_net_1 ), .Y(
        N_282));
    DFN1E1 \acqtime[9]  (.D(noisedata[9]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[9]_net_1 ));
    OAI1 \CS_RNO_0[6]  (.A(\CS[6]_net_1 ), .B(timer_top_0_clk_en_noise)
        , .C(top_code_0_noise_rst_0), .Y(\CS_srsts_i_0[6] ));
    OA1 \CS_i_0_RNO[0]  (.A(\CS_li[0] ), .B(timer_top_0_clk_en_noise), 
        .C(top_code_0_noise_rst), .Y(\CS_i_0_RNO_0[0] ));
    DFN1 state_over_n (.D(state_over_n_RNO_1), .CLK(GLA), .Q(
        noisestate_0_state_over_n));
    NOR2A \CS_RNO[1]  (.A(top_code_0_noise_rst_0), .B(
        \CS_srsts_i_0[1] ), .Y(\CS_RNO_2[1] ));
    MX2 \timecount_1_RNO[3]  (.A(N_64), .B(N_243), .S(N_280), .Y(
        \timecount_5[3] ));
    VCC VCC_i (.Y(VCC));
    DFN1E1 \timecount_1[7]  (.D(\timecount_5[7] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[7]));
    DFN1E1 \dectime[12]  (.D(noisedata[12]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[12]_net_1 ));
    OAI1 \CS_RNO_0[2]  (.A(\CS[2]_net_1 ), .B(timer_top_0_clk_en_noise)
        , .C(top_code_0_noise_rst_0), .Y(\CS_srsts_i_0[2] ));
    DFN1E1 \acqtime[2]  (.D(noisedata[2]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[2]_net_1 ));
    NOR2 \timecount_1_RNO[12]  (.A(N_280), .B(N_73), .Y(
        \timecount_5[12] ));
    MX2B rt_sw_RNO_0 (.A(noisestate_0_rt_sw), .B(\CS[5]_net_1 ), .S(
        N_300), .Y(N_114));
    DFN1 dumpon_ctr (.D(dumpon_ctr_RNO_0_net_1), .CLK(GLA), .Q(
        noisestate_0_dumpon_ctr));
    NOR2 \CS_RNID768[6]  (.A(\CS[7]_net_1 ), .B(\CS[6]_net_1 ), .Y(
        N_302));
    DFN1E1 \timecount_1[15]  (.D(\timecount_5[15] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[15]));
    NOR2A \CS_RNO_1[5]  (.A(timer_top_0_clk_en_noise), .B(
        \CS[4]_net_1 ), .Y(N_295));
    DFN1E1 \dectime[6]  (.D(noisedata[6]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[6]_net_1 ));
    DFN1 dumpoff_ctr (.D(dumpoff_ctr_RNO_2), .CLK(GLA), .Q(
        noisestate_0_dumpoff_ctr));
    MX2C \timecount_1_RNO_0[1]  (.A(\acqtime[1]_net_1 ), .B(
        \dectime[1]_net_1 ), .S(N_245), .Y(N_62));
    MX2C \timecount_1_RNO_0[13]  (.A(\dectime[13]_net_1 ), .B(
        \acqtime[13]_net_1 ), .S(\CS[4]_net_1 ), .Y(N_74));
    MX2 \timecount_1_RNO_0[11]  (.A(\acqtime[11]_net_1 ), .B(
        \dectime[11]_net_1 ), .S(N_245), .Y(N_72));
    MX2C \timecount_1_RNO[0]  (.A(N_61), .B(top_code_0_noise_rst), .S(
        N_280), .Y(\timecount_5[0] ));
    DFN1E1 \timecount_1[6]  (.D(\timecount_5[6] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[6]));
    DFN1 n_acq (.D(n_acq_RNO_net_1), .CLK(GLA), .Q(noisestate_0_n_acq));
    OR2A \CS_RNIT5UE[6]  (.A(top_code_0_noise_rst), .B(N_302), .Y(
        un1_dumpoff_ctr_2_sqmuxa));
    NOR2B \CS_RNI1CQA_0[1]  (.A(top_code_0_noise_rst), .B(
        \CS[1]_net_1 ), .Y(N_243));
    NOR2 sw_acq2_RNO_1 (.A(\CS[4]_net_1 ), .B(\CS[3]_net_1 ), .Y(N_286)
        );
    DFN1 \CS[7]  (.D(\CS_RNO_2[7] ), .CLK(GLA), .Q(\CS[7]_net_1 ));
    NOR2 \timecount_1_RNO[15]  (.A(N_280), .B(N_76), .Y(
        \timecount_5[15] ));
    DFN1 \CS[6]  (.D(\CS_RNO_2[6] ), .CLK(GLA), .Q(\CS[6]_net_1 ));
    DFN1E1 \dectime[0]  (.D(noisedata[0]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[0]_net_1 ));
    AO1B state_over_n_RNO (.A(noisestate_0_state_over_n), .B(N_302), 
        .C(top_code_0_noise_rst_0), .Y(state_over_n_RNO_1));
    MX2C \timecount_1_RNO_0[0]  (.A(\acqtime[0]_net_1 ), .B(
        \dectime[0]_net_1 ), .S(N_245), .Y(N_61));
    DFN1E1 \acqtime[1]  (.D(noisedata[1]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[1]_net_1 ));
    MX2C \timecount_1_RNO_0[6]  (.A(\acqtime[6]_net_1 ), .B(
        \dectime[6]_net_1 ), .S(N_245), .Y(N_67));
    OA1C \CS_RNO[2]  (.A(timer_top_0_clk_en_noise), .B(\CS[1]_net_1 ), 
        .C(\CS_srsts_i_0[2] ), .Y(\CS_RNO_2[2] ));
    GND GND_i_0 (.Y(GND_0));
    MX2C \timecount_1_RNO_0[8]  (.A(\dectime[8]_net_1 ), .B(
        \acqtime[8]_net_1 ), .S(\CS[4]_net_1 ), .Y(N_69));
    DFN1E1 \acqtime[0]  (.D(noisedata[0]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[0]_net_1 ));
    NOR2 \timecount_1_RNO[1]  (.A(N_280), .B(N_62), .Y(
        \timecount_5[1] ));
    OR3B \CS_i_0_RNI028F[0]  (.A(\CS_li[0] ), .B(
        top_code_0_noise_rst_0), .C(\CS[5]_net_1 ), .Y(
        \timecount_cnst[4] ));
    MX2 sw_acq2_RNO_0 (.A(noisestate_0_sw_acq2), .B(N_286), .S(N_300), 
        .Y(N_112));
    AO1 dumpoff_ctr_RNO_0 (.A(noisestate_0_dumpoff_ctr), .B(N_302), .C(
        \CS[5]_net_1 ), .Y(N_116));
    DFN1E1 \acqtime[8]  (.D(noisedata[8]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[8]_net_1 ));
    DFN1 \CS[2]  (.D(\CS_RNO_2[2] ), .CLK(GLA), .Q(\CS[2]_net_1 ));
    DFN1E1 \dectime[11]  (.D(noisedata[11]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[11]_net_1 ));
    DFN1E1 \dectime[4]  (.D(noisedata[4]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[4]_net_1 ));
    NOR2 \timecount_1_RNO[13]  (.A(N_280), .B(N_74), .Y(
        \timecount_5[13] ));
    DFN1E1 \acqtime[5]  (.D(noisedata[5]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[5]_net_1 ));
    AO1A n_acq_RNO_0 (.A(\CS[5]_net_1 ), .B(noisestate_0_n_acq), .C(
        \CS[4]_net_1 ), .Y(N_133));
    DFN1E1 \timecount_1[9]  (.D(\timecount_5[9] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[9]));
    OR2B \CS_RNI4OQA[4]  (.A(top_code_0_noise_rst), .B(\CS[4]_net_1 ), 
        .Y(N_245));
    DFN1E1 \dectime[3]  (.D(noisedata[3]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[3]_net_1 ));
    NOR2 \timecount_1_RNO[14]  (.A(N_280), .B(N_75), .Y(
        \timecount_5[14] ));
    OAI1 \CS_RNIM9TE[2]  (.A(\CS[2]_net_1 ), .B(\CS[4]_net_1 ), .C(
        top_code_0_noise_rst), .Y(N_280));
    DFN1 \CS[5]  (.D(\CS_RNO_2[5] ), .CLK(GLA), .Q(\CS[5]_net_1 ));
    MX2C \timecount_1_RNO[2]  (.A(N_63), .B(\timecount_cnst[2] ), .S(
        N_280), .Y(\timecount_5[2] ));
    OAI1 \CS_RNO_0[3]  (.A(\CS[3]_net_1 ), .B(timer_top_0_clk_en_noise)
        , .C(top_code_0_noise_rst_0), .Y(\CS_srsts_i_0[3] ));
    DFN1E1 \acqtime[3]  (.D(noisedata[3]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[3]_net_1 ));
    DFN1E1 \timecount_1[3]  (.D(\timecount_5[3] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[3]));
    NOR2B n_acq_RNO (.A(top_code_0_noise_rst), .B(N_133), .Y(
        n_acq_RNO_net_1));
    MX2 \timecount_1_RNO[9]  (.A(N_70), .B(N_243), .S(N_280), .Y(
        \timecount_5[9] ));
    DFN1 rt_sw (.D(rt_sw_RNO_2), .CLK(GLA), .Q(noisestate_0_rt_sw));
    DFN1E1 \dectime[14]  (.D(noisedata[14]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[14]_net_1 ));
    DFN1E1 \dectime[7]  (.D(noisedata[7]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[7]_net_1 ));
    OA1C \CS_RNO[6]  (.A(timer_top_0_clk_en_noise), .B(\CS[5]_net_1 ), 
        .C(\CS_srsts_i_0[6] ), .Y(\CS_RNO_2[6] ));
    MX2 \timecount_1_RNO[11]  (.A(N_72), .B(N_243), .S(N_280), .Y(
        \timecount_5[11] ));
    MX2C \timecount_1_RNO_0[7]  (.A(\acqtime[7]_net_1 ), .B(
        \dectime[7]_net_1 ), .S(N_245), .Y(N_68));
    MX2C \timecount_1_RNO[8]  (.A(N_69), .B(\timecount_cnst[4] ), .S(
        N_280), .Y(\timecount_5[8] ));
    DFN1E1 \dectime[9]  (.D(noisedata[9]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[9]_net_1 ));
    DFN1E1 \acqtime[13]  (.D(noisedata[13]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[13]_net_1 ));
    DFN1E1 \acqtime[12]  (.D(noisedata[12]), .CLK(GLA), .E(
        acqtime_1_sqmuxa_net_1), .Q(\acqtime[12]_net_1 ));
    DFN1E1 \timecount_1[4]  (.D(\timecount_5[4] ), .CLK(GLA), .E(
        un1_dumpoff_ctr_2_sqmuxa), .Q(timecount_1[4]));
    DFN1E1 \dectime[5]  (.D(noisedata[5]), .CLK(GLA), .E(
        acqtime_0_sqmuxa_net_1), .Q(\dectime[5]_net_1 ));
    MX2C \timecount_1_RNO_0[15]  (.A(\acqtime[15]_net_1 ), .B(
        \dectime[15]_net_1 ), .S(N_245), .Y(N_76));
    NOR2A acqtime_1_sqmuxa (.A(top_code_0_nstateload), .B(
        top_code_0_nstatechoice), .Y(acqtime_1_sqmuxa_net_1));
    MX2C \timecount_1_RNO_0[14]  (.A(\acqtime[14]_net_1 ), .B(
        \dectime[14]_net_1 ), .S(N_245), .Y(N_75));
    
endmodule


module dds_change(
       un1_top_code_0_3_0,
       GLA,
       top_code_0_pluse_rst,
       net_45,
       net_33_0,
       plusestate_0_dds_config,
       scalestate_0_dds_conf,
       scanstate_0_dds_conf,
       net_27,
       dds_change_0_dds_conf,
       un1_change_2,
       dds_change_0_dds_rst
    );
input  [1:0] un1_top_code_0_3_0;
input  GLA;
input  top_code_0_pluse_rst;
input  net_45;
input  net_33_0;
input  plusestate_0_dds_config;
input  scalestate_0_dds_conf;
input  scanstate_0_dds_conf;
input  net_27;
output dds_change_0_dds_conf;
output un1_change_2;
output dds_change_0_dds_rst;

    wire dds_rst_6, ddsrstin3_m, ddsrstin2_m, ddsrstin1_m, dds_conf_6, 
        dds_confin3_m, dds_confin2_m, dds_confin1_m, N_5, N_6, 
        dds_conf_RNO_net_1, dds_rst_RNO_net_1, GND, VCC, GND_0, VCC_0;
    
    OR3A dds_rst_RNO_4 (.A(net_33_0), .B(un1_top_code_0_3_0[0]), .C(
        un1_top_code_0_3_0[1]), .Y(ddsrstin1_m));
    GND GND_i_0 (.Y(GND_0));
    MX2 dds_conf_RNO_0 (.A(dds_change_0_dds_conf), .B(dds_conf_6), .S(
        un1_change_2), .Y(N_6));
    OR2B dds_rst_RNO_3 (.A(un1_top_code_0_3_0[0]), .B(net_45), .Y(
        ddsrstin2_m));
    VCC VCC_i (.Y(VCC));
    OR3C dds_rst_RNO_1 (.A(ddsrstin3_m), .B(ddsrstin2_m), .C(
        ddsrstin1_m), .Y(dds_rst_6));
    NOR2B dds_rst_RNO (.A(net_27), .B(N_5), .Y(dds_rst_RNO_net_1));
    OR3A dds_conf_RNO_4 (.A(scanstate_0_dds_conf), .B(
        un1_top_code_0_3_0[0]), .C(un1_top_code_0_3_0[1]), .Y(
        dds_confin1_m));
    GND GND_i (.Y(GND));
    VCC VCC_i_0 (.Y(VCC_0));
    OR2B dds_rst_RNO_2 (.A(un1_top_code_0_3_0[1]), .B(
        top_code_0_pluse_rst), .Y(ddsrstin3_m));
    DFN1 dds_conf (.D(dds_conf_RNO_net_1), .CLK(GLA), .Q(
        dds_change_0_dds_conf));
    OR2B dds_conf_RNO_2 (.A(un1_top_code_0_3_0[1]), .B(
        plusestate_0_dds_config), .Y(dds_confin3_m));
    OR3C dds_conf_RNO_1 (.A(dds_confin3_m), .B(dds_confin2_m), .C(
        dds_confin1_m), .Y(dds_conf_6));
    OR2B un1_change_2_inst_1 (.A(un1_top_code_0_3_0[1]), .B(
        un1_top_code_0_3_0[0]), .Y(un1_change_2));
    DFN1 dds_rst (.D(dds_rst_RNO_net_1), .CLK(GLA), .Q(
        dds_change_0_dds_rst));
    NOR2B dds_conf_RNO (.A(net_27), .B(N_6), .Y(dds_conf_RNO_net_1));
    MX2 dds_rst_RNO_0 (.A(dds_change_0_dds_rst), .B(dds_rst_6), .S(
        un1_change_2), .Y(N_5));
    OR2B dds_conf_RNO_3 (.A(un1_top_code_0_3_0[0]), .B(
        scalestate_0_dds_conf), .Y(dds_confin2_m));
    
endmodule


module NMR_TOP(
       zcs2,
       xwe,
       ddsfqud,
       ddsreset,
       ddswclk,
       cal_out,
       ddsdata,
       OCX40MHz,
       ddsclkout,
       interupt,
       rt_sw,
       soft_dump,
       sw_acq1,
       sw_acq2,
       dumpon,
       dumpoff,
       Q1Q8,
       Q3Q6,
       Q4Q5,
       Q2Q7,
       calcuinter,
       tri_ctrl,
       sigtimeup,
       k1,
       k2,
       gpio,
       pulse_start,
       pd_pulse_en,
       XRD,
       Acq_clk,
       sd_acq_en,
       s_acq180,
       GLA,
       xa,
       xd,
       relayclose_on,
       ADC
    );
input  zcs2;
input  xwe;
output ddsfqud;
output ddsreset;
output ddswclk;
output cal_out;
output ddsdata;
input  OCX40MHz;
input  ddsclkout;
output interupt;
output rt_sw;
output soft_dump;
output sw_acq1;
output sw_acq2;
output dumpon;
output dumpoff;
output Q1Q8;
output Q3Q6;
output Q4Q5;
output Q2Q7;
output calcuinter;
input  tri_ctrl;
output sigtimeup;
output k1;
output k2;
input  gpio;
output pulse_start;
output pd_pulse_en;
input  XRD;
output Acq_clk;
output sd_acq_en;
output s_acq180;
output GLA;
input  [18:0] xa;
inout  [15:0] xd;
output [15:0] relayclose_on;
input  [11:0] ADC;

    wire net_27, top_code_0_pluse_noise_ctrl, noisestate_0_n_acq, 
        plusestate_0_pluse_acq, n_acq_change_0_n_acq_start, 
        top_code_0_noise_rst, top_code_0_pluse_rst, 
        n_acq_change_0_n_rst_n, timer_top_0_clk_en_pluse, 
        plusestate_0_soft_d, plusestate_0_sw_acq1, \timecount_1_1[0] , 
        \timecount_1_1[1] , \timecount_1_1[2] , \timecount_1_1[3] , 
        \timecount_1_1[4] , \timecount_1_1[5] , \timecount_1_1[6] , 
        \timecount_1_1[7] , \timecount_1_1[8] , \timecount_1_1[9] , 
        \timecount_1_1[10] , \timecount_1_1[11] , \timecount_1_1[12] , 
        \timecount_1_1[13] , \timecount_1_1[14] , \timecount_1_1[15] , 
        plusestate_0_off_test, \plusedata[0] , \plusedata[1] , 
        \plusedata[2] , \plusedata[3] , \plusedata[4] , \plusedata[5] , 
        \plusedata[6] , \plusedata[7] , \plusedata[8] , \plusedata[9] , 
        \plusedata[10] , \plusedata[11] , \plusedata[12] , 
        \plusedata[13] , \plusedata[14] , \plusedata[15] , 
        top_code_0_pluseload, top_code_0_pluse_lc, 
        plusestate_0_state_over_n, plusestate_0_dds_config, 
        plusestate_0_tetw_pluse, \change[0] , \change[1] , 
        dds_change_0_dds_rst, net_33, net_45, dds_change_0_dds_conf, 
        scalestate_0_dds_conf, bri_dump_sw_0_reset_out, 
        bri_dump_sw_0_phase_ctr, net_51, top_code_0_bridge_load, 
        \bri_datain[0] , \bri_datain[1] , \bri_datain[2] , 
        \bri_datain[3] , \bri_datain[4] , \bri_datain[5] , 
        \bri_datain[6] , \bri_datain[7] , \bri_datain[8] , 
        \bri_datain[9] , \bri_datain[10] , \bri_datain[11] , 
        \bri_datain[12] , \bri_datain[13] , \bri_datain[14] , 
        \bri_datain[15] , \halfdata[0] , \halfdata[1] , \halfdata[2] , 
        \halfdata[3] , \halfdata[4] , \halfdata[5] , \halfdata[6] , 
        \halfdata[7] , top_code_0_dds_load, top_code_0_dds_choice, 
        \dds_configdata[0] , \dds_configdata[1] , \dds_configdata[2] , 
        \dds_configdata[3] , \dds_configdata[4] , \dds_configdata[5] , 
        \dds_configdata[6] , \dds_configdata[7] , \dds_configdata[8] , 
        \dds_configdata[9] , \dds_configdata[10] , 
        \dds_configdata[11] , \dds_configdata[12] , 
        \dds_configdata[13] , \dds_configdata[14] , 
        \dds_configdata[15] , Signal_Noise_Acq_0_acq_clk, 
        top_code_0_acqclken, GPMI_0_code_en, top_code_0_scan_start, 
        top_code_0_noise_start, top_code_0_cal_load, \cal_data[0] , 
        \cal_data[1] , \cal_data[2] , \cal_data[3] , \cal_data[4] , 
        \cal_data[5] , \s_acqnum_0[0] , \s_acqnum_0[1] , 
        \s_acqnum_0[2] , \s_acqnum_0[3] , \s_acqnum_0[4] , 
        \s_acqnum_0[5] , \s_acqnum_0[6] , \s_acqnum_0[7] , 
        \s_acqnum_0[8] , \s_acqnum_0[9] , \s_acqnum_0[10] , 
        \s_acqnum_0[11] , \s_acqnum_0[12] , \s_acqnum_0[13] , 
        \s_acqnum_0[14] , \s_acqnum_0[15] , top_code_0_s_load, 
        top_code_0_scale_rst, top_code_0_scale_start, 
        top_code_0_scaleload, top_code_0_pn_change, 
        top_code_0_dumpload, \scaledatain[0] , \scaledatain[1] , 
        \scaledatain[2] , \scaledatain[3] , \scaledatain[4] , 
        \scaledatain[5] , \scaledatain[6] , \scaledatain[7] , 
        \scaledatain[8] , \scaledatain[9] , \scaledatain[10] , 
        \scaledatain[11] , \scaledatain[12] , \scaledatain[13] , 
        \scaledatain[14] , \scaledatain[15] , \scalechoice[0] , 
        \scalechoice[1] , \scalechoice[2] , \scalechoice[3] , 
        \scalechoice[4] , \dump_cho[0] , \dump_cho[1] , \dump_cho[2] , 
        \dumpdata[0] , \dumpdata[1] , \dumpdata[2] , \dumpdata[3] , 
        \dumpdata[4] , \dumpdata[5] , \dumpdata[6] , \dumpdata[7] , 
        \dumpdata[8] , \dumpdata[9] , \dumpdata[10] , \dumpdata[11] , 
        \scaleddsdiv[0] , \scaleddsdiv[1] , \scaleddsdiv[2] , 
        \scaleddsdiv[3] , \scaleddsdiv[4] , \scaleddsdiv[5] , 
        top_code_0_pluse_scale, top_code_0_pluse_str, \sigtimedata[0] , 
        \sigtimedata[1] , \sigtimedata[2] , \sigtimedata[3] , 
        \sigtimedata[4] , \sigtimedata[5] , \sigtimedata[6] , 
        \sigtimedata[7] , \sigtimedata[8] , \sigtimedata[9] , 
        \sigtimedata[10] , \sigtimedata[11] , \sigtimedata[12] , 
        \sigtimedata[13] , \sigtimedata[14] , \sigtimedata[15] , 
        top_code_0_sigrst, top_code_0_scanchoice, top_code_0_scanload, 
        \scandata[0] , \scandata[1] , \scandata[2] , \scandata[3] , 
        \scandata[4] , \scandata[5] , \scandata[6] , \scandata[7] , 
        \scandata[8] , \scandata[9] , \scandata[10] , \scandata[11] , 
        \scandata[12] , \scandata[13] , \scandata[14] , \scandata[15] , 
        top_code_0_nstateload, top_code_0_nstatechoice, \noisedata[0] , 
        \noisedata[1] , \noisedata[2] , \noisedata[3] , \noisedata[4] , 
        \noisedata[5] , \noisedata[6] , \noisedata[7] , \noisedata[8] , 
        \noisedata[9] , \noisedata[10] , \noisedata[11] , 
        \noisedata[12] , \noisedata[13] , \noisedata[14] , 
        \noisedata[15] , top_code_0_state_1ms_rst_n, 
        top_code_0_state_1ms_start, \state_1ms_lc[0] , 
        \state_1ms_lc[1] , \state_1ms_lc[2] , \state_1ms_lc[3] , 
        top_code_0_state_1ms_load, \state_1ms_data[0] , 
        \state_1ms_data[1] , \state_1ms_data[2] , \state_1ms_data[3] , 
        \state_1ms_data[4] , \state_1ms_data[5] , \state_1ms_data[6] , 
        \state_1ms_data[7] , \state_1ms_data[8] , \state_1ms_data[9] , 
        \state_1ms_data[10] , \state_1ms_data[11] , 
        \state_1ms_data[12] , \state_1ms_data[13] , 
        \state_1ms_data[14] , \state_1ms_data[15] , top_code_0_n_load, 
        top_code_0_n_s_ctrl, \n_divnum[0] , \n_divnum[1] , 
        \n_divnum[2] , \n_divnum[3] , \n_divnum[4] , \n_divnum[5] , 
        \n_divnum[6] , \n_divnum[7] , \n_divnum[8] , \n_divnum[9] , 
        \s_periodnum[0] , \s_periodnum[1] , \s_periodnum[2] , 
        \s_periodnum[3] , \n_acqnum[0] , \n_acqnum[1] , \n_acqnum[2] , 
        \n_acqnum[3] , \n_acqnum[4] , \n_acqnum[5] , \n_acqnum[6] , 
        \n_acqnum[7] , \n_acqnum[8] , \n_acqnum[9] , \n_acqnum[10] , 
        \n_acqnum[11] , \sd_sacq_choice[0] , \sd_sacq_choice[1] , 
        \sd_sacq_choice[2] , \sd_sacq_choice[3] , \sd_sacq_data[0] , 
        \sd_sacq_data[1] , \sd_sacq_data[2] , \sd_sacq_data[3] , 
        \sd_sacq_data[4] , \sd_sacq_data[5] , \sd_sacq_data[6] , 
        \sd_sacq_data[7] , \sd_sacq_data[8] , \sd_sacq_data[9] , 
        \sd_sacq_data[10] , \sd_sacq_data[11] , \sd_sacq_data[12] , 
        \sd_sacq_data[13] , \sd_sacq_data[14] , \sd_sacq_data[15] , 
        top_code_0_sd_sacq_load, \pd_pluse_choice[0] , 
        \pd_pluse_choice[1] , \pd_pluse_choice[2] , 
        \pd_pluse_choice[3] , top_code_0_pd_pluse_load, 
        \pd_pluse_data[0] , \pd_pluse_data[1] , \pd_pluse_data[2] , 
        \pd_pluse_data[3] , \pd_pluse_data[4] , \pd_pluse_data[5] , 
        \pd_pluse_data[6] , \pd_pluse_data[7] , \pd_pluse_data[8] , 
        \pd_pluse_data[9] , \pd_pluse_data[10] , \pd_pluse_data[11] , 
        \pd_pluse_data[12] , \pd_pluse_data[13] , \pd_pluse_data[14] , 
        \pd_pluse_data[15] , top_code_0_RAM_Rd_rst, top_code_0_n_rd_en, 
        \s_addchoice[0] , \s_addchoice[1] , \s_addchoice[2] , 
        \s_addchoice[3] , \s_addchoice[4] , top_code_0_dump_sustain, 
        scalestate_0_dump_sustain_ctrl, AND2_1_Y, 
        dump_sustain_timer_0_start, clk_5K, scanstate_0_soft_d, 
        scanstate_0_rt_sw, scanstate_0_sw_acq2, 
        scanstate_0_state_over_n, scanstate_0_dds_conf, 
        scanstate_0_dumpoff_ctr, noisestate_0_soft_d, 
        noisestate_0_rt_sw, noisestate_0_sw_acq2, 
        noisestate_0_state_over_n, noisestate_0_dumpon_ctr, 
        noisestate_0_dumpoff_ctr, nsctrl_choice_0_soft_d, 
        nsctrl_choice_0_rt_sw, nsctrl_choice_0_sw_acq2, 
        nsctrl_choice_0_intertodsp, nsctrl_choice_0_dumpon_ctr, 
        nsctrl_choice_0_dumpoff_ctr, nsctrl_choice_0_dumponoff_rst, 
        bri_div_start_0, state_1ms_0_pluse_start, 
        bri_dump_sw_0_off_test, state1ms_choice_0_dump_start, 
        state_1ms_0_dump_start, bri_dump_sw_0_dump_start, 
        state1ms_choice_0_reset_out, state_1ms_0_reset_out, 
        state1ms_choice_0_bri_cycle, state_1ms_0_bri_cycle, 
        state_1ms_0_rt_sw, rt_sw_net_1, state_1ms_0_soft_dump, 
        soft_dump_net_1, bri_dump_sw_0_dumpoff_ctr, scalestate_0_s_acq, 
        scalestate_0_long_opentime, timer_top_0_clk_en_scan, 
        timer_top_0_clk_en_st1ms, timer_top_0_clk_en_scale, 
        timer_top_0_clk_en_noise, \timecount_0[0] , \timecount_0[1] , 
        \timecount_0[2] , \timecount_0[3] , \timecount_0[4] , 
        \timecount_0[5] , \timecount_0[6] , \timecount_0[7] , 
        \timecount_0[8] , \timecount_0[9] , \timecount_0[10] , 
        \timecount_0[11] , \timecount_0[12] , \timecount_0[13] , 
        \timecount_0[14] , \timecount_0[15] , \timecount_0[16] , 
        \timecount_0[17] , \timecount_0[18] , \timecount_0[19] , 
        \timecount[0] , \timecount[1] , \timecount[2] , \timecount[3] , 
        \timecount[4] , \timecount[5] , \timecount[6] , \timecount[7] , 
        \timecount[8] , \timecount[9] , \timecount[10] , 
        \timecount[11] , \timecount[12] , \timecount[13] , 
        \timecount[14] , \timecount[15] , \timecount[16] , 
        \timecount[17] , \timecount[18] , \timecount[19] , 
        \timecount[20] , \timecount[21] , \timecount_1_0[0] , 
        \timecount_1_0[1] , \timecount_1_0[2] , \timecount_1_0[3] , 
        \timecount_1_0[4] , \timecount_1_0[5] , \timecount_1_0[6] , 
        \timecount_1_0[7] , \timecount_1_0[8] , \timecount_1_0[9] , 
        \timecount_1_0[10] , \timecount_1_0[11] , \timecount_1_0[12] , 
        \timecount_1_0[13] , \timecount_1_0[14] , \timecount_1_0[15] , 
        \timecount_1[0] , \timecount_1[1] , \timecount_1[2] , 
        \timecount_1[3] , \timecount_1[4] , \timecount_1[5] , 
        \timecount_1[6] , \timecount_1[7] , \timecount_1[8] , 
        \timecount_1[9] , \timecount_1[10] , \timecount_1[11] , 
        \timecount_1[12] , \timecount_1[13] , \timecount_1[14] , 
        \timecount_1[15] , scalestate_0_tetw_pluse, 
        scalestate_0_pluse_start, scalestate_0_off_test, 
        scalestate_0_dump_start, scalestate_0_pn_out, 
        scalestate_0_dumpoff_ctr, bri_dump_sw_0_tetw_pluse, 
        scan_scale_sw_0_s_start, scanstate_0_s_acq, 
        s_acq_change_0_s_load, scalestate_0_load_out, 
        s_acq_change_0_s_rst, \s_acqnum[0] , \s_acqnum[1] , 
        \s_acqnum[2] , \s_acqnum[3] , \s_acqnum[4] , \s_acqnum[5] , 
        \s_acqnum[6] , \s_acqnum[7] , \s_acqnum[8] , \s_acqnum[9] , 
        \s_acqnum[10] , \s_acqnum[11] , \s_acqnum[12] , \s_acqnum[13] , 
        \s_acqnum[14] , \s_acqnum[15] , \s_acqnum_1[0] , 
        \s_acqnum_1[1] , \s_acqnum_1[2] , \s_acqnum_1[3] , 
        \s_acqnum_1[4] , \s_acqnum_1[5] , \s_acqnum_1[6] , 
        \s_acqnum_1[7] , \s_acqnum_1[8] , \s_acqnum_1[9] , 
        \s_acqnum_1[10] , \s_acqnum_1[11] , \s_stripnum[0] , 
        \s_stripnum[1] , \s_stripnum[2] , \s_stripnum[3] , 
        \s_stripnum[4] , \s_stripnum[5] , \s_stripnum[6] , 
        \s_stripnum[7] , \s_stripnum[8] , \s_stripnum[9] , 
        \s_stripnum[10] , \s_stripnum[11] , \strippluse[0] , 
        \strippluse[1] , \strippluse[2] , \strippluse[3] , 
        \strippluse[4] , \strippluse[5] , \strippluse[6] , 
        \strippluse[7] , \strippluse[8] , \strippluse[9] , 
        \strippluse[10] , \strippluse[11] , scanstate_0_calctrl, 
        OR2_1_Y, OR2_2_Y, scalestate_0_rt_sw, scalestate_0_soft_d, 
        scalestate_0_sw_acq1, scalestate_0_sw_acq2, \dataout_0[12] , 
        \dataout_0[13] , \dataout_0[14] , \dataout_0[15] , VCC, GND, 
        \GPMI_0.tri_state_0.xd_1 , \dataout_0[3] , \dataout_0[4] , 
        \dataout_0[9] , \dataout_0[10] , \dataout_0[0] , 
        \dataout_0[2] , \dataout_0[6] , \dataout_0[8] , \dataout_0[1] , 
        \dataout_0[5] , \dataout_0[7] , \dataout_0[11] , 
        DUMP_0_dump_off, DUMP_0_dump_on, DUMP_OFF_1_dump_off, 
        DUMP_ON_0_dump_on, \i_0_0[1] , \i_4[1] , DUMP_OFF_0_dump_off, 
        \xd_in[0] , \xd_in[1] , \xd_in[2] , \xd_in[3] , \xd_in[4] , 
        \xd_in[5] , \xd_in[6] , \xd_in[7] , \xd_in[8] , \xd_in[9] , 
        \xd_in[10] , \xd_in[11] , \xd_in[12] , \xd_in[13] , 
        \xd_in[14] , \xd_in[15] , zcs2_c, xwe_c, ddsfqud_c, ddsreset_c, 
        ddswclk_c, cal_out_c, ddsdata_c, OCX40MHz_c, ddsclkout_c, 
        interupt_c, rt_sw_c, soft_dump_c, sw_acq1_c, sw_acq2_c, 
        dumpon_c, dumpoff_c, Q1Q8_c, Q3Q6_c, Q4Q5_c, Q2Q7_c, 
        calcuinter_c, tri_ctrl_c, sigtimeup_c, k1_c, k2_c, gpio_c, 
        pulse_start_c, pd_pulse_en_c, XRD_c, Acq_clk_c, sd_acq_en_c, 
        s_acq180_c, GLA_net_1, \xa_c[0] , \xa_c[1] , \xa_c[2] , 
        \xa_c[3] , \xa_c[4] , \xa_c[5] , \xa_c[6] , \xa_c[7] , 
        \xa_c[8] , \xa_c[9] , \xa_c[10] , \xa_c[11] , \xa_c[12] , 
        \xa_c[13] , \xa_c[14] , \xa_c[15] , \xa_c[16] , \xa_c[17] , 
        \xa_c[18] , \relayclose_on_c[0] , \relayclose_on_c[1] , 
        \relayclose_on_c[2] , \relayclose_on_c[3] , 
        \relayclose_on_c[4] , \relayclose_on_c[5] , 
        \relayclose_on_c[6] , \relayclose_on_c[7] , 
        \relayclose_on_c[8] , \relayclose_on_c[9] , 
        \relayclose_on_c[10] , \relayclose_on_c[11] , 
        \relayclose_on_c[12] , \relayclose_on_c[13] , 
        \relayclose_on_c[14] , \relayclose_on_c[15] , \ADC_c[0] , 
        \ADC_c[1] , \ADC_c[2] , \ADC_c[3] , \ADC_c[4] , \ADC_c[5] , 
        \ADC_c[6] , \ADC_c[7] , \ADC_c[8] , \ADC_c[9] , \ADC_c[10] , 
        \ADC_c[11] , \un1_GPMI_0_1[0] , \un1_GPMI_0_1[1] , 
        \un1_GPMI_0_1[2] , \un1_GPMI_0_1[3] , \un1_GPMI_0_1[4] , 
        \un1_GPMI_0_1[5] , \un1_GPMI_0_1[6] , \un1_GPMI_0_1[7] , 
        \un1_GPMI_0_1[8] , \un1_GPMI_0_1[9] , \un1_GPMI_0_1[10] , 
        \un1_GPMI_0_1[11] , \un1_GPMI_0_1[13] , \un1_GPMI_0_1[14] , 
        \un1_GPMI_0_1[15] , \un1_GPMI_0_1[12] , clk_4f_en, 
        \dds_change_0.un1_change_2 , PLUSE_0_bri_cycle, 
        \un1_GPMI_0_1_0[2] , \un1_GPMI_0_1_0[1] , \un1_GPMI_0_1_0[0] , 
        \xa_c_0[7] , \xa_c_0[0] , s_acq_change_0_s_load_0, 
        timer_top_0_clk_en_scale_0, top_code_0_n_s_ctrl_0, 
        top_code_0_n_s_ctrl_1, top_code_0_state_1ms_rst_n_0, 
        top_code_0_bridge_load_0, bri_dump_sw_0_reset_out_0, net_33_0, 
        \un1_top_code_0_3_0[1] , \un1_top_code_0_3_0[0] , 
        n_acq_change_0_n_rst_n_0, top_code_0_pluse_rst_0, 
        top_code_0_noise_rst_0, GND_0, VCC_0;
    
    OUTBUF Q4Q5_pad (.D(Q4Q5_c), .PAD(Q4Q5));
    NOR2A \xd_pad_RNISLFD[14]  (.A(\xd_in[14] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[14] ));
    NOR2A \xd_pad_RNIE8Q8[7]  (.A(\xd_in[7] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[7] ));
    NOR2A \xd_pad_RNI78Q8_0[0]  (.A(\xd_in[0] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[0] ));
    INBUF \ADC_pad[0]  (.PAD(ADC[0]), .Y(\ADC_c[0] ));
    state1ms_choice state1ms_choice_0 (.state1ms_choice_0_bri_cycle(
        state1ms_choice_0_bri_cycle), .state1ms_choice_0_dump_start(
        state1ms_choice_0_dump_start), .bri_div_start_0(
        bri_div_start_0), .state1ms_choice_0_reset_out(
        state1ms_choice_0_reset_out), .rt_sw_c(rt_sw_c), .GLA(
        GLA_net_1), .soft_dump_c(soft_dump_c), .state_1ms_0_soft_dump(
        state_1ms_0_soft_dump), .soft_dump_net_1(soft_dump_net_1), 
        .state_1ms_0_rt_sw(state_1ms_0_rt_sw), .rt_sw_net_1(
        rt_sw_net_1), .state_1ms_0_reset_out(state_1ms_0_reset_out), 
        .bri_dump_sw_0_reset_out_0(bri_dump_sw_0_reset_out_0), 
        .state_1ms_0_pluse_start(state_1ms_0_pluse_start), 
        .bri_dump_sw_0_off_test(bri_dump_sw_0_off_test), 
        .state_1ms_0_dump_start(state_1ms_0_dump_start), 
        .bri_dump_sw_0_dump_start(bri_dump_sw_0_dump_start), 
        .top_code_0_state_1ms_start(top_code_0_state_1ms_start), 
        .state_1ms_0_bri_cycle(state_1ms_0_bri_cycle), 
        .PLUSE_0_bri_cycle(PLUSE_0_bri_cycle), .net_27(net_27));
    top_code top_code_0 (.plusedata({\plusedata[15] , \plusedata[14] , 
        \plusedata[13] , \plusedata[12] , \plusedata[11] , 
        \plusedata[10] , \plusedata[9] , \plusedata[8] , 
        \plusedata[7] , \plusedata[6] , \plusedata[5] , \plusedata[4] , 
        \plusedata[3] , \plusedata[2] , \plusedata[1] , \plusedata[0] })
        , .s_acqnum_0({\s_acqnum_0[15] , \s_acqnum_0[14] , 
        \s_acqnum_0[13] , \s_acqnum_0[12] , \s_acqnum_0[11] , 
        \s_acqnum_0[10] , \s_acqnum_0[9] , \s_acqnum_0[8] , 
        \s_acqnum_0[7] , \s_acqnum_0[6] , \s_acqnum_0[5] , 
        \s_acqnum_0[4] , \s_acqnum_0[3] , \s_acqnum_0[2] , 
        \s_acqnum_0[1] , \s_acqnum_0[0] }), .s_addchoice({
        \s_addchoice[4] , \s_addchoice[3] , \s_addchoice[2] , 
        \s_addchoice[1] , \s_addchoice[0] }), .s_periodnum({
        \s_periodnum[3] , \s_periodnum[2] , \s_periodnum[1] , 
        \s_periodnum[0] }), .scalechoice({\scalechoice[4] , 
        \scalechoice[3] , \scalechoice[2] , \scalechoice[1] , 
        \scalechoice[0] }), .scaledatain({\scaledatain[15] , 
        \scaledatain[14] , \scaledatain[13] , \scaledatain[12] , 
        \scaledatain[11] , \scaledatain[10] , \scaledatain[9] , 
        \scaledatain[8] , \scaledatain[7] , \scaledatain[6] , 
        \scaledatain[5] , \scaledatain[4] , \scaledatain[3] , 
        \scaledatain[2] , \scaledatain[1] , \scaledatain[0] }), 
        .scaleddsdiv({\scaleddsdiv[5] , \scaleddsdiv[4] , 
        \scaleddsdiv[3] , \scaleddsdiv[2] , \scaleddsdiv[1] , 
        \scaleddsdiv[0] }), .scandata({\scandata[15] , \scandata[14] , 
        \scandata[13] , \scandata[12] , \scandata[11] , \scandata[10] , 
        \scandata[9] , \scandata[8] , \scandata[7] , \scandata[6] , 
        \scandata[5] , \scandata[4] , \scandata[3] , \scandata[2] , 
        \scandata[1] , \scandata[0] }), .sd_sacq_choice({
        \sd_sacq_choice[3] , \sd_sacq_choice[2] , \sd_sacq_choice[1] , 
        \sd_sacq_choice[0] }), .sd_sacq_data({\sd_sacq_data[15] , 
        \sd_sacq_data[14] , \sd_sacq_data[13] , \sd_sacq_data[12] , 
        \sd_sacq_data[11] , \sd_sacq_data[10] , \sd_sacq_data[9] , 
        \sd_sacq_data[8] , \sd_sacq_data[7] , \sd_sacq_data[6] , 
        \sd_sacq_data[5] , \sd_sacq_data[4] , \sd_sacq_data[3] , 
        \sd_sacq_data[2] , \sd_sacq_data[1] , \sd_sacq_data[0] }), 
        .sigtimedata({\sigtimedata[15] , \sigtimedata[14] , 
        \sigtimedata[13] , \sigtimedata[12] , \sigtimedata[11] , 
        \sigtimedata[10] , \sigtimedata[9] , \sigtimedata[8] , 
        \sigtimedata[7] , \sigtimedata[6] , \sigtimedata[5] , 
        \sigtimedata[4] , \sigtimedata[3] , \sigtimedata[2] , 
        \sigtimedata[1] , \sigtimedata[0] }), .state_1ms_data({
        \state_1ms_data[15] , \state_1ms_data[14] , 
        \state_1ms_data[13] , \state_1ms_data[12] , 
        \state_1ms_data[11] , \state_1ms_data[10] , 
        \state_1ms_data[9] , \state_1ms_data[8] , \state_1ms_data[7] , 
        \state_1ms_data[6] , \state_1ms_data[5] , \state_1ms_data[4] , 
        \state_1ms_data[3] , \state_1ms_data[2] , \state_1ms_data[1] , 
        \state_1ms_data[0] }), .state_1ms_lc({\state_1ms_lc[3] , 
        \state_1ms_lc[2] , \state_1ms_lc[1] , \state_1ms_lc[0] }), 
        .bri_datain({\bri_datain[15] , \bri_datain[14] , 
        \bri_datain[13] , \bri_datain[12] , \bri_datain[11] , 
        \bri_datain[10] , \bri_datain[9] , \bri_datain[8] , 
        \bri_datain[7] , \bri_datain[6] , \bri_datain[5] , 
        \bri_datain[4] , \bri_datain[3] , \bri_datain[2] , 
        \bri_datain[1] , \bri_datain[0] }), .cal_data({\cal_data[5] , 
        \cal_data[4] , \cal_data[3] , \cal_data[2] , \cal_data[1] , 
        \cal_data[0] }), .change({\change[1] , \change[0] }), 
        .dds_configdata({\dds_configdata[15] , \dds_configdata[14] , 
        \dds_configdata[13] , \dds_configdata[12] , 
        \dds_configdata[11] , \dds_configdata[10] , 
        \dds_configdata[9] , \dds_configdata[8] , \dds_configdata[7] , 
        \dds_configdata[6] , \dds_configdata[5] , \dds_configdata[4] , 
        \dds_configdata[3] , \dds_configdata[2] , \dds_configdata[1] , 
        \dds_configdata[0] }), .dump_cho({\dump_cho[2] , \dump_cho[1] , 
        \dump_cho[0] }), .dumpdata({\dumpdata[11] , \dumpdata[10] , 
        \dumpdata[9] , \dumpdata[8] , \dumpdata[7] , \dumpdata[6] , 
        \dumpdata[5] , \dumpdata[4] , \dumpdata[3] , \dumpdata[2] , 
        \dumpdata[1] , \dumpdata[0] }), .halfdata({\halfdata[7] , 
        \halfdata[6] , \halfdata[5] , \halfdata[4] , \halfdata[3] , 
        \halfdata[2] , \halfdata[1] , \halfdata[0] }), .n_acqnum({
        \n_acqnum[11] , \n_acqnum[10] , \n_acqnum[9] , \n_acqnum[8] , 
        \n_acqnum[7] , \n_acqnum[6] , \n_acqnum[5] , \n_acqnum[4] , 
        \n_acqnum[3] , \n_acqnum[2] , \n_acqnum[1] , \n_acqnum[0] }), 
        .n_divnum({\n_divnum[9] , \n_divnum[8] , \n_divnum[7] , 
        \n_divnum[6] , \n_divnum[5] , \n_divnum[4] , \n_divnum[3] , 
        \n_divnum[2] , \n_divnum[1] , \n_divnum[0] }), .noisedata({
        \noisedata[15] , \noisedata[14] , \noisedata[13] , 
        \noisedata[12] , \noisedata[11] , \noisedata[10] , 
        \noisedata[9] , \noisedata[8] , \noisedata[7] , \noisedata[6] , 
        \noisedata[5] , \noisedata[4] , \noisedata[3] , \noisedata[2] , 
        \noisedata[1] , \noisedata[0] }), .pd_pluse_choice({
        \pd_pluse_choice[3] , \pd_pluse_choice[2] , 
        \pd_pluse_choice[1] , \pd_pluse_choice[0] }), .pd_pluse_data({
        \pd_pluse_data[15] , \pd_pluse_data[14] , \pd_pluse_data[13] , 
        \pd_pluse_data[12] , \pd_pluse_data[11] , \pd_pluse_data[10] , 
        \pd_pluse_data[9] , \pd_pluse_data[8] , \pd_pluse_data[7] , 
        \pd_pluse_data[6] , \pd_pluse_data[5] , \pd_pluse_data[4] , 
        \pd_pluse_data[3] , \pd_pluse_data[2] , \pd_pluse_data[1] , 
        \pd_pluse_data[0] }), .un1_GPMI_0_1({\un1_GPMI_0_1[15] , 
        \un1_GPMI_0_1[14] , \un1_GPMI_0_1[13] , \un1_GPMI_0_1[12] , 
        \un1_GPMI_0_1[11] , \un1_GPMI_0_1[10] , \un1_GPMI_0_1[9] , 
        \un1_GPMI_0_1[8] , \un1_GPMI_0_1[7] , \un1_GPMI_0_1[6] , 
        \un1_GPMI_0_1[5] , \un1_GPMI_0_1[4] , \un1_GPMI_0_1[3] , 
        \un1_GPMI_0_1[2] , \un1_GPMI_0_1[1] , \un1_GPMI_0_1[0] }), 
        .relayclose_on_c({\relayclose_on_c[15] , \relayclose_on_c[14] , 
        \relayclose_on_c[13] , \relayclose_on_c[12] , 
        \relayclose_on_c[11] , \relayclose_on_c[10] , 
        \relayclose_on_c[9] , \relayclose_on_c[8] , 
        \relayclose_on_c[7] , \relayclose_on_c[6] , 
        \relayclose_on_c[5] , \relayclose_on_c[4] , 
        \relayclose_on_c[3] , \relayclose_on_c[2] , 
        \relayclose_on_c[1] , \relayclose_on_c[0] }), .xa_c_0_0(
        \xa_c_0[0] ), .xa_c_0_7(\xa_c_0[7] ), .xa_c({\xa_c[18] , 
        \xa_c[17] , \xa_c[16] , \xa_c[15] , \xa_c[14] , \xa_c[13] , 
        \xa_c[12] , \xa_c[11] , \xa_c[10] , \xa_c[9] , \xa_c[8] , 
        \xa_c[7] , \xa_c[6] , \xa_c[5] , \xa_c[4] , \xa_c[3] , 
        \xa_c[2] , \xa_c[1] , \xa_c[0] }), .un1_GPMI_0_1_0({
        \un1_GPMI_0_1_0[2] , \un1_GPMI_0_1_0[1] , \un1_GPMI_0_1_0[0] })
        , .un1_top_code_0_3_0({\un1_top_code_0_3_0[1] , 
        \un1_top_code_0_3_0[0] }), .net_33(net_33), 
        .top_code_0_noise_rst(top_code_0_noise_rst), 
        .top_code_0_bridge_load(top_code_0_bridge_load), 
        .top_code_0_scale_start(top_code_0_scale_start), 
        .top_code_0_pn_change(top_code_0_pn_change), 
        .top_code_0_scanload(top_code_0_scanload), 
        .top_code_0_acqclken(top_code_0_acqclken), 
        .top_code_0_state_1ms_rst_n(top_code_0_state_1ms_rst_n), 
        .top_code_0_scaleload(top_code_0_scaleload), 
        .top_code_0_scan_start(top_code_0_scan_start), 
        .top_code_0_n_load(top_code_0_n_load), .top_code_0_n_rd_en(
        top_code_0_n_rd_en), .top_code_0_n_s_ctrl(top_code_0_n_s_ctrl), 
        .top_code_0_RAM_Rd_rst(top_code_0_RAM_Rd_rst), 
        .top_code_0_noise_start(top_code_0_noise_start), 
        .top_code_0_dds_choice(top_code_0_dds_choice), 
        .top_code_0_dumpload(top_code_0_dumpload), 
        .top_code_0_pluseload(top_code_0_pluseload), 
        .top_code_0_scanchoice(top_code_0_scanchoice), 
        .top_code_0_pluse_scale(top_code_0_pluse_scale), 
        .top_code_0_state_1ms_load(top_code_0_state_1ms_load), 
        .top_code_0_sd_sacq_load(top_code_0_sd_sacq_load), 
        .top_code_0_pd_pluse_load(top_code_0_pd_pluse_load), 
        .top_code_0_nstateload(top_code_0_nstateload), 
        .top_code_0_pluse_lc(top_code_0_pluse_lc), .top_code_0_sigrst(
        top_code_0_sigrst), .top_code_0_s_load(top_code_0_s_load), 
        .top_code_0_cal_load(top_code_0_cal_load), 
        .top_code_0_nstatechoice(top_code_0_nstatechoice), 
        .top_code_0_pluse_noise_ctrl(top_code_0_pluse_noise_ctrl), 
        .top_code_0_dump_sustain(top_code_0_dump_sustain), .k1_c(k1_c), 
        .k2_c(k2_c), .top_code_0_pluse_rst(top_code_0_pluse_rst), 
        .top_code_0_pluse_str(top_code_0_pluse_str), 
        .top_code_0_state_1ms_start(top_code_0_state_1ms_start), 
        .GPMI_0_code_en(GPMI_0_code_en), .top_code_0_scale_rst(
        top_code_0_scale_rst), .top_code_0_dds_load(
        top_code_0_dds_load), .top_code_0_n_s_ctrl_0(
        top_code_0_n_s_ctrl_0), .top_code_0_n_s_ctrl_1(
        top_code_0_n_s_ctrl_1), .top_code_0_state_1ms_rst_n_0(
        top_code_0_state_1ms_rst_n_0), .net_27(net_27), 
        .top_code_0_bridge_load_0(top_code_0_bridge_load_0), .net_33_0(
        net_33_0), .top_code_0_pluse_rst_0(top_code_0_pluse_rst_0), 
        .GLA(GLA_net_1), .top_code_0_noise_rst_0(
        top_code_0_noise_rst_0));
    BIBUF \xd_pad[11]  (.PAD(xd[11]), .D(\dataout_0[11] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[11] ));
    INBUF \xa_pad[4]  (.PAD(xa[4]), .Y(\xa_c[4] ));
    OR2 OR2_2 (.A(nsctrl_choice_0_dumponoff_rst), .B(
        scalestate_0_dump_sustain_ctrl), .Y(OR2_2_Y));
    INBUF xwe_pad (.PAD(xwe), .Y(xwe_c));
    scan_scale_sw scan_scale_sw_0 (.change({\change[1] }), 
        .un1_top_code_0_3_0({\un1_top_code_0_3_0[0] }), .ddsclkout_c(
        ddsclkout_c), .net_27(net_27), .scan_scale_sw_0_s_start(
        scan_scale_sw_0_s_start), .sd_acq_en_c(sd_acq_en_c), 
        .scanstate_0_s_acq(scanstate_0_s_acq));
    NOR2A \xd_pad_RNIB8Q8[4]  (.A(\xd_in[4] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[4] ));
    INBUF \xa_pad[14]  (.PAD(xa[14]), .Y(\xa_c[14] ));
    OUTBUF Q2Q7_pad (.D(Q2Q7_c), .PAD(Q2Q7));
    OUTBUF calcuinter_pad (.D(calcuinter_c), .PAD(calcuinter));
    OUTBUF dumpon_pad (.D(dumpon_c), .PAD(dumpon));
    AND2 AND2_1 (.A(scalestate_0_dump_sustain_ctrl), .B(
        top_code_0_dump_sustain), .Y(AND2_1_Y));
    OUTBUF k2_pad (.D(k2_c), .PAD(k2));
    DDS DDS_0 (.dds_configdata({\dds_configdata[15] , 
        \dds_configdata[14] , \dds_configdata[13] , 
        \dds_configdata[12] , \dds_configdata[11] , 
        \dds_configdata[10] , \dds_configdata[9] , \dds_configdata[8] , 
        \dds_configdata[7] , \dds_configdata[6] , \dds_configdata[5] , 
        \dds_configdata[4] , \dds_configdata[3] , \dds_configdata[2] , 
        \dds_configdata[1] , \dds_configdata[0] }), 
        .top_code_0_dds_load(top_code_0_dds_load), 
        .top_code_0_dds_choice(top_code_0_dds_choice), .ddswclk_c(
        ddswclk_c), .ddsfqud_c(ddsfqud_c), .ddsdata_c(ddsdata_c), 
        .ddsreset_c(ddsreset_c), .dds_change_0_dds_conf(
        dds_change_0_dds_conf), .dds_change_0_dds_rst(
        dds_change_0_dds_rst), .GLA(GLA_net_1));
    INBUF zcs2_pad (.PAD(zcs2), .Y(zcs2_c));
    BIBUF \xd_pad[7]  (.PAD(xd[7]), .D(\dataout_0[7] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[7] ));
    timer_top timer_top_0 (.timecount_1_0({\timecount_1_0[15] , 
        \timecount_1_0[14] , \timecount_1_0[13] , \timecount_1_0[12] , 
        \timecount_1_0[11] , \timecount_1_0[10] , \timecount_1_0[9] , 
        \timecount_1_0[8] , \timecount_1_0[7] , \timecount_1_0[6] , 
        \timecount_1_0[5] , \timecount_1_0[4] , \timecount_1_0[3] , 
        \timecount_1_0[2] , \timecount_1_0[1] , \timecount_1_0[0] }), 
        .timecount_1_1({\timecount_1_1[15] , \timecount_1_1[14] , 
        \timecount_1_1[13] , \timecount_1_1[12] , \timecount_1_1[11] , 
        \timecount_1_1[10] , \timecount_1_1[9] , \timecount_1_1[8] , 
        \timecount_1_1[7] , \timecount_1_1[6] , \timecount_1_1[5] , 
        \timecount_1_1[4] , \timecount_1_1[3] , \timecount_1_1[2] , 
        \timecount_1_1[1] , \timecount_1_1[0] }), .timecount({
        \timecount[21] , \timecount[20] , \timecount[19] , 
        \timecount[18] , \timecount[17] , \timecount[16] , 
        \timecount[15] , \timecount[14] , \timecount[13] , 
        \timecount[12] , \timecount[11] , \timecount[10] , 
        \timecount[9] , \timecount[8] , \timecount[7] , \timecount[6] , 
        \timecount[5] , \timecount[4] , \timecount[3] , \timecount[2] , 
        \timecount[1] , \timecount[0] }), .timecount_0({
        \timecount_0[19] , \timecount_0[18] , \timecount_0[17] , 
        \timecount_0[16] , \timecount_0[15] , \timecount_0[14] , 
        \timecount_0[13] , \timecount_0[12] , \timecount_0[11] , 
        \timecount_0[10] , \timecount_0[9] , \timecount_0[8] , 
        \timecount_0[7] , \timecount_0[6] , \timecount_0[5] , 
        \timecount_0[4] , \timecount_0[3] , \timecount_0[2] , 
        \timecount_0[1] , \timecount_0[0] }), .timecount_1({
        \timecount_1[15] , \timecount_1[14] , \timecount_1[13] , 
        \timecount_1[12] , \timecount_1[11] , \timecount_1[10] , 
        \timecount_1[9] , \timecount_1[8] , \timecount_1[7] , 
        \timecount_1[6] , \timecount_1[5] , \timecount_1[4] , 
        \timecount_1[3] , \timecount_1[2] , \timecount_1[1] , 
        \timecount_1[0] }), .timer_top_0_clk_en_scale_0(
        timer_top_0_clk_en_scale_0), .plusestate_0_state_over_n(
        plusestate_0_state_over_n), .top_code_0_scan_start(
        top_code_0_scan_start), .top_code_0_noise_start(
        top_code_0_noise_start), .top_code_0_scale_start(
        top_code_0_scale_start), .top_code_0_state_1ms_start(
        top_code_0_state_1ms_start), .scanstate_0_state_over_n(
        scanstate_0_state_over_n), .noisestate_0_state_over_n(
        noisestate_0_state_over_n), .scalestate_0_tetw_pluse(
        scalestate_0_tetw_pluse), .top_code_0_pluse_str(
        top_code_0_pluse_str), .timer_top_0_clk_en_st1ms(
        timer_top_0_clk_en_st1ms), .timer_top_0_clk_en_scan(
        timer_top_0_clk_en_scan), .timer_top_0_clk_en_scale(
        timer_top_0_clk_en_scale), .timer_top_0_clk_en_pluse(
        timer_top_0_clk_en_pluse), .timer_top_0_clk_en_noise(
        timer_top_0_clk_en_noise), .net_27(net_27), .GLA(GLA_net_1));
    OUTBUF Acq_clk_pad (.D(Acq_clk_c), .PAD(Acq_clk));
    NOR2A \xd_pad_RNIO5FD[10]  (.A(\xd_in[10] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[10] ));
    INBUF gpio_pad (.PAD(gpio), .Y(gpio_c));
    OUTBUF ddsfqud_pad (.D(ddsfqud_c), .PAD(ddsfqud));
    OUTBUF ddsdata_pad (.D(ddsdata_c), .PAD(ddsdata));
    BIBUF \xd_pad[4]  (.PAD(xd[4]), .D(\dataout_0[4] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[4] ));
    NOR2A \xd_pad_RNID8Q8[6]  (.A(\xd_in[6] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[6] ));
    OUTBUF \relayclose_on_pad[10]  (.D(\relayclose_on_c[10] ), .PAD(
        relayclose_on[10]));
    INBUF \xa_pad[16]  (.PAD(xa[16]), .Y(\xa_c[16] ));
    NOR2A \xd_pad_RNIF8Q8[8]  (.A(\xd_in[8] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[8] ));
    OR2 OR2_0 (.A(DUMP_0_dump_on), .B(DUMP_ON_0_dump_on), .Y(dumpon_c));
    OUTBUF interupt_pad (.D(interupt_c), .PAD(interupt));
    Signal_Noise_Acq Signal_Noise_Acq_0 (.dataout_0({\dataout_0[15] , 
        \dataout_0[14] , \dataout_0[13] , \dataout_0[12] , 
        \dataout_0[11] , \dataout_0[10] , \dataout_0[9] , 
        \dataout_0[8] , \dataout_0[7] , \dataout_0[6] , \dataout_0[5] , 
        \dataout_0[4] , \dataout_0[3] , \dataout_0[2] , \dataout_0[1] , 
        \dataout_0[0] }), .n_divnum({\n_divnum[9] , \n_divnum[8] , 
        \n_divnum[7] , \n_divnum[6] , \n_divnum[5] , \n_divnum[4] , 
        \n_divnum[3] , \n_divnum[2] , \n_divnum[1] , \n_divnum[0] }), 
        .n_acqnum({\n_acqnum[11] , \n_acqnum[10] , \n_acqnum[9] , 
        \n_acqnum[8] , \n_acqnum[7] , \n_acqnum[6] , \n_acqnum[5] , 
        \n_acqnum[4] , \n_acqnum[3] , \n_acqnum[2] , \n_acqnum[1] , 
        \n_acqnum[0] }), .s_addchoice({\s_addchoice[4] , 
        \s_addchoice[3] , \s_addchoice[2] , \s_addchoice[1] , 
        \s_addchoice[0] }), .s_acqnum({\s_acqnum[15] , \s_acqnum[14] , 
        \s_acqnum[13] , \s_acqnum[12] , \s_acqnum[11] , \s_acqnum[10] , 
        \s_acqnum[9] , \s_acqnum[8] , \s_acqnum[7] , \s_acqnum[6] , 
        \s_acqnum[5] , \s_acqnum[4] , \s_acqnum[3] , \s_acqnum[2] , 
        \s_acqnum[1] , \s_acqnum[0] }), .s_periodnum({\s_periodnum[3] , 
        \s_periodnum[2] , \s_periodnum[1] , \s_periodnum[0] }), 
        .s_stripnum({\s_stripnum[11] , \s_stripnum[10] , 
        \s_stripnum[9] , \s_stripnum[8] , \s_stripnum[7] , 
        \s_stripnum[6] , \s_stripnum[5] , \s_stripnum[4] , 
        \s_stripnum[3] , \s_stripnum[2] , \s_stripnum[1] , 
        \s_stripnum[0] }), .ADC_c({\ADC_c[11] , \ADC_c[10] , 
        \ADC_c[9] , \ADC_c[8] , \ADC_c[7] , \ADC_c[6] , \ADC_c[5] , 
        \ADC_c[4] , \ADC_c[3] , \ADC_c[2] , \ADC_c[1] , \ADC_c[0] }), 
        .Signal_Noise_Acq_0_acq_clk(Signal_Noise_Acq_0_acq_clk), 
        .XRD_c(XRD_c), .n_acq_change_0_n_rst_n_0(
        n_acq_change_0_n_rst_n_0), .top_code_0_n_rd_en(
        top_code_0_n_rd_en), .n_acq_change_0_n_rst_n(
        n_acq_change_0_n_rst_n), .top_code_0_n_load(top_code_0_n_load), 
        .n_acq_change_0_n_acq_start(n_acq_change_0_n_acq_start), 
        .Signal_Noise_Acq_VCC(VCC), .Signal_Noise_Acq_GND(GND), 
        .top_code_0_RAM_Rd_rst(top_code_0_RAM_Rd_rst), 
        .s_acq_change_0_s_rst(s_acq_change_0_s_rst), .ddsclkout_c(
        ddsclkout_c), .scan_scale_sw_0_s_start(scan_scale_sw_0_s_start)
        , .s_acq_change_0_s_load_0(s_acq_change_0_s_load_0), 
        .s_acq_change_0_s_load(s_acq_change_0_s_load), .GLA(GLA_net_1), 
        .top_code_0_n_s_ctrl(top_code_0_n_s_ctrl), 
        .top_code_0_n_s_ctrl_1(top_code_0_n_s_ctrl_1), 
        .top_code_0_n_s_ctrl_0(top_code_0_n_s_ctrl_0));
    NOR2A \xd_pad_RNIRHFD[13]  (.A(\xd_in[13] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[13] ));
    OUTBUF \relayclose_on_pad[2]  (.D(\relayclose_on_c[2] ), .PAD(
        relayclose_on[2]));
    GND GND_i (.Y(GND));
    OUTBUF \relayclose_on_pad[14]  (.D(\relayclose_on_c[14] ), .PAD(
        relayclose_on[14]));
    VCC VCC_i_0 (.Y(VCC_0));
    INBUF XRD_pad (.PAD(XRD), .Y(XRD_c));
    bri_dump_sw bri_dump_sw_0 (.bri_dump_sw_0_dump_start(
        bri_dump_sw_0_dump_start), .bri_dump_sw_0_dumpoff_ctr(
        bri_dump_sw_0_dumpoff_ctr), .bri_dump_sw_0_off_test(
        bri_dump_sw_0_off_test), .bri_dump_sw_0_phase_ctr(
        bri_dump_sw_0_phase_ctr), .pulse_start_c(pulse_start_c), 
        .bri_dump_sw_0_reset_out(bri_dump_sw_0_reset_out), 
        .bri_dump_sw_0_tetw_pluse(bri_dump_sw_0_tetw_pluse), .net_45(
        net_45), .top_code_0_pluse_rst(top_code_0_pluse_rst), 
        .scalestate_0_tetw_pluse(scalestate_0_tetw_pluse), 
        .scalestate_0_pluse_start(scalestate_0_pluse_start), 
        .scalestate_0_pn_out(scalestate_0_pn_out), 
        .top_code_0_pn_change(top_code_0_pn_change), 
        .scalestate_0_off_test(scalestate_0_off_test), 
        .plusestate_0_off_test(plusestate_0_off_test), 
        .scalestate_0_dumpoff_ctr(scalestate_0_dumpoff_ctr), 
        .plusestate_0_tetw_pluse(plusestate_0_tetw_pluse), 
        .top_code_0_pluse_scale(top_code_0_pluse_scale), 
        .scalestate_0_dump_start(scalestate_0_dump_start), 
        .plusestate_0_soft_d(plusestate_0_soft_d), .net_27(net_27), 
        .GLA(GLA_net_1), .bri_dump_sw_0_reset_out_0(
        bri_dump_sw_0_reset_out_0));
    INBUF \ADC_pad[3]  (.PAD(ADC[3]), .Y(\ADC_c[3] ));
    INBUF \xa_pad[5]  (.PAD(xa[5]), .Y(\xa_c[5] ));
    INBUF \ADC_pad[9]  (.PAD(ADC[9]), .Y(\ADC_c[9] ));
    INBUF \xa_pad[10]  (.PAD(xa[10]), .Y(\xa_c[10] ));
    OUTBUF \relayclose_on_pad[11]  (.D(\relayclose_on_c[11] ), .PAD(
        relayclose_on[11]));
    BIBUF \xd_pad[2]  (.PAD(xd[2]), .D(\dataout_0[2] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[2] ));
    INBUF \xa_pad[18]  (.PAD(xa[18]), .Y(\xa_c[18] ));
    OUTBUF \relayclose_on_pad[7]  (.D(\relayclose_on_c[7] ), .PAD(
        relayclose_on[7]));
    BIBUF \xd_pad[13]  (.PAD(xd[13]), .D(\dataout_0[13] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[13] ));
    dump_sustain_timer dump_sustain_timer_0 (
        .dump_sustain_timer_0_start(dump_sustain_timer_0_start), 
        .clk_5K(clk_5K), .AND2_1_Y(AND2_1_Y), 
        .scalestate_0_dump_sustain_ctrl(scalestate_0_dump_sustain_ctrl)
        );
    INBUF tri_ctrl_pad (.PAD(tri_ctrl), .Y(tri_ctrl_c));
    OUTBUF \relayclose_on_pad[4]  (.D(\relayclose_on_c[4] ), .PAD(
        relayclose_on[4]));
    NOR2A \xd_pad_RNI78Q8[0]  (.A(\xd_in[0] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1_0[0] ));
    INBUF \xa_pad[15]  (.PAD(xa[15]), .Y(\xa_c[15] ));
    INBUF \xa_pad[17]  (.PAD(xa[17]), .Y(\xa_c[17] ));
    CAL CAL_0 (.cal_data({\cal_data[5] , \cal_data[4] , \cal_data[3] , 
        \cal_data[2] , \cal_data[1] , \cal_data[0] }), 
        .scanstate_0_calctrl(scanstate_0_calctrl), .net_33(net_33), 
        .cal_out_c(cal_out_c), .ddsclkout_c(ddsclkout_c), .GLA(
        GLA_net_1), .top_code_0_cal_load(top_code_0_cal_load));
    OUTBUF k1_pad (.D(k1_c), .PAD(k1));
    OUTBUF dumpoff_pad (.D(dumpoff_c), .PAD(dumpoff));
    OUTBUF \relayclose_on_pad[13]  (.D(\relayclose_on_c[13] ), .PAD(
        relayclose_on[13]));
    VCC VCC_i (.Y(VCC));
    INBUF \ADC_pad[1]  (.PAD(ADC[1]), .Y(\ADC_c[1] ));
    PLUSE PLUSE_0 (.bri_datain({\bri_datain[15] , \bri_datain[14] , 
        \bri_datain[13] , \bri_datain[12] , \bri_datain[11] , 
        \bri_datain[10] , \bri_datain[9] , \bri_datain[8] , 
        \bri_datain[7] , \bri_datain[6] , \bri_datain[5] , 
        \bri_datain[4] , \bri_datain[3] , \bri_datain[2] , 
        \bri_datain[1] , \bri_datain[0] }), .halfdata({\halfdata[7] , 
        \halfdata[6] , \halfdata[5] , \halfdata[4] , \halfdata[3] , 
        \halfdata[2] , \halfdata[1] , \halfdata[0] }), 
        .top_code_0_bridge_load(top_code_0_bridge_load), 
        .top_code_0_bridge_load_0(top_code_0_bridge_load_0), .Q4Q5_c(
        Q4Q5_c), .Q2Q7_c(Q2Q7_c), .PLUSE_0_bri_cycle(PLUSE_0_bri_cycle)
        , .bri_dump_sw_0_phase_ctr(bri_dump_sw_0_phase_ctr), .net_51(
        net_51), .clk_4f_en(clk_4f_en), .pulse_start_c(pulse_start_c), 
        .ddsclkout_c(ddsclkout_c), .bri_dump_sw_0_reset_out(
        bri_dump_sw_0_reset_out), .bri_dump_sw_0_reset_out_0(
        bri_dump_sw_0_reset_out_0), .Q3Q6_c(Q3Q6_c), .Q1Q8_c(Q1Q8_c), 
        .GLA(GLA_net_1));
    BIBUF \xd_pad[12]  (.PAD(xd[12]), .D(\dataout_0[12] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[12] ));
    state_1ms state_1ms_0 (.state_1ms_data({\state_1ms_data[15] , 
        \state_1ms_data[14] , \state_1ms_data[13] , 
        \state_1ms_data[12] , \state_1ms_data[11] , 
        \state_1ms_data[10] , \state_1ms_data[9] , \state_1ms_data[8] , 
        \state_1ms_data[7] , \state_1ms_data[6] , \state_1ms_data[5] , 
        \state_1ms_data[4] , \state_1ms_data[3] , \state_1ms_data[2] , 
        \state_1ms_data[1] , \state_1ms_data[0] }), .timecount_0({
        \timecount_0[19] , \timecount_0[18] , \timecount_0[17] , 
        \timecount_0[16] , \timecount_0[15] , \timecount_0[14] , 
        \timecount_0[13] , \timecount_0[12] , \timecount_0[11] , 
        \timecount_0[10] , \timecount_0[9] , \timecount_0[8] , 
        \timecount_0[7] , \timecount_0[6] , \timecount_0[5] , 
        \timecount_0[4] , \timecount_0[3] , \timecount_0[2] , 
        \timecount_0[1] , \timecount_0[0] }), .state_1ms_lc({
        \state_1ms_lc[3] , \state_1ms_lc[2] , \state_1ms_lc[1] , 
        \state_1ms_lc[0] }), .GLA(GLA_net_1), .state_1ms_0_reset_out(
        state_1ms_0_reset_out), .top_code_0_state_1ms_rst_n(
        top_code_0_state_1ms_rst_n), .top_code_0_state_1ms_load(
        top_code_0_state_1ms_load), .state_1ms_0_bri_cycle(
        state_1ms_0_bri_cycle), .state_1ms_0_pluse_start(
        state_1ms_0_pluse_start), .state_1ms_0_rt_sw(state_1ms_0_rt_sw)
        , .state_1ms_0_soft_dump(state_1ms_0_soft_dump), 
        .state_1ms_0_dump_start(state_1ms_0_dump_start), 
        .top_code_0_state_1ms_rst_n_0(top_code_0_state_1ms_rst_n_0), 
        .timer_top_0_clk_en_st1ms(timer_top_0_clk_en_st1ms));
    sd_acq_top sd_acq_top_0 (.sd_sacq_choice({\sd_sacq_choice[3] , 
        \sd_sacq_choice[2] , \sd_sacq_choice[1] , \sd_sacq_choice[0] })
        , .sd_sacq_data({\sd_sacq_data[15] , \sd_sacq_data[14] , 
        \sd_sacq_data[13] , \sd_sacq_data[12] , \sd_sacq_data[11] , 
        \sd_sacq_data[10] , \sd_sacq_data[9] , \sd_sacq_data[8] , 
        \sd_sacq_data[7] , \sd_sacq_data[6] , \sd_sacq_data[5] , 
        \sd_sacq_data[4] , \sd_sacq_data[3] , \sd_sacq_data[2] , 
        \sd_sacq_data[1] , \sd_sacq_data[0] }), .i_4_1(\i_4[1] ), 
        .i_0_0({\i_0_0[1] }), .sd_acq_en_c(sd_acq_en_c), .net_27(
        net_27), .scalestate_0_s_acq(scalestate_0_s_acq), 
        .top_code_0_sd_sacq_load(top_code_0_sd_sacq_load), .s_acq180_c(
        s_acq180_c), .scalestate_0_long_opentime(
        scalestate_0_long_opentime), .GLA(GLA_net_1), .ddsclkout_c(
        ddsclkout_c));
    INBUF OCX40MHz_pad (.PAD(OCX40MHz), .Y(OCX40MHz_c));
    BIBUF \xd_pad[5]  (.PAD(xd[5]), .D(\dataout_0[5] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[5] ));
    CLKBUF ddsclkout_pad (.PAD(ddsclkout), .Y(ddsclkout_c));
    INBUF \xa_pad[8]  (.PAD(xa[8]), .Y(\xa_c[8] ));
    OUTBUF sigtimeup_pad (.D(sigtimeup_c), .PAD(sigtimeup));
    INBUF \ADC_pad[5]  (.PAD(ADC[5]), .Y(\ADC_c[5] ));
    OUTBUF \relayclose_on_pad[8]  (.D(\relayclose_on_c[8] ), .PAD(
        relayclose_on[8]));
    DUMP_OFF_DUMP_OFF_0_1 DUMP_OFF_1 (.nsctrl_choice_0_dumpoff_ctr(
        nsctrl_choice_0_dumpoff_ctr), .nsctrl_choice_0_dumponoff_rst(
        nsctrl_choice_0_dumponoff_rst), .DUMP_OFF_1_dump_off(
        DUMP_OFF_1_dump_off), .GLA(GLA_net_1));
    OUTBUF sw_acq2_pad (.D(sw_acq2_c), .PAD(sw_acq2));
    INBUF \ADC_pad[10]  (.PAD(ADC[10]), .Y(\ADC_c[10] ));
    INBUF \xa_pad[11]  (.PAD(xa[11]), .Y(\xa_c[11] ));
    INBUF \ADC_pad[8]  (.PAD(ADC[8]), .Y(\ADC_c[8] ));
    BIBUF \xd_pad[8]  (.PAD(xd[8]), .D(\dataout_0[8] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[8] ));
    OUTBUF \relayclose_on_pad[0]  (.D(\relayclose_on_c[0] ), .PAD(
        relayclose_on[0]));
    OUTBUF GLA_pad (.D(GLA_net_1), .PAD(GLA));
    OUTBUF rt_sw_pad (.D(rt_sw_c), .PAD(rt_sw));
    INBUF \xa_pad[7]  (.PAD(xa[7]), .Y(\xa_c[7] ));
    INBUF \xa_pad[6]  (.PAD(xa[6]), .Y(\xa_c[6] ));
    BIBUF \xd_pad[6]  (.PAD(xd[6]), .D(\dataout_0[6] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[6] ));
    OUTBUF \relayclose_on_pad[9]  (.D(\relayclose_on_c[9] ), .PAD(
        relayclose_on[9]));
    BIBUF \xd_pad[9]  (.PAD(xd[9]), .D(\dataout_0[9] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[9] ));
    scalestate scalestate_0 (.timecount({\timecount[21] , 
        \timecount[20] , \timecount[19] , \timecount[18] , 
        \timecount[17] , \timecount[16] , \timecount[15] , 
        \timecount[14] , \timecount[13] , \timecount[12] , 
        \timecount[11] , \timecount[10] , \timecount[9] , 
        \timecount[8] , \timecount[7] , \timecount[6] , \timecount[5] , 
        \timecount[4] , \timecount[3] , \timecount[2] , \timecount[1] , 
        \timecount[0] }), .scaledatain({\scaledatain[15] , 
        \scaledatain[14] , \scaledatain[13] , \scaledatain[12] , 
        \scaledatain[11] , \scaledatain[10] , \scaledatain[9] , 
        \scaledatain[8] , \scaledatain[7] , \scaledatain[6] , 
        \scaledatain[5] , \scaledatain[4] , \scaledatain[3] , 
        \scaledatain[2] , \scaledatain[1] , \scaledatain[0] }), 
        .strippluse({\strippluse[11] , \strippluse[10] , 
        \strippluse[9] , \strippluse[8] , \strippluse[7] , 
        \strippluse[6] , \strippluse[5] , \strippluse[4] , 
        \strippluse[3] , \strippluse[2] , \strippluse[1] , 
        \strippluse[0] }), .s_acqnum_1({\s_acqnum_1[11] , 
        \s_acqnum_1[10] , \s_acqnum_1[9] , \s_acqnum_1[8] , 
        \s_acqnum_1[7] , \s_acqnum_1[6] , \s_acqnum_1[5] , 
        \s_acqnum_1[4] , \s_acqnum_1[3] , \s_acqnum_1[2] , 
        \s_acqnum_1[1] , \s_acqnum_1[0] }), .scalechoice({
        \scalechoice[4] , \scalechoice[3] , \scalechoice[2] , 
        \scalechoice[1] , \scalechoice[0] }), .net_45(net_45), 
        .timer_top_0_clk_en_scale(timer_top_0_clk_en_scale), 
        .scalestate_0_dump_start(scalestate_0_dump_start), 
        .scalestate_0_soft_d(scalestate_0_soft_d), .scalestate_0_rt_sw(
        scalestate_0_rt_sw), .net_51(net_51), 
        .scalestate_0_long_opentime(scalestate_0_long_opentime), 
        .scalestate_0_s_acq(scalestate_0_s_acq), 
        .scalestate_0_pluse_start(scalestate_0_pluse_start), 
        .s_acq180_c(s_acq180_c), .scalestate_0_tetw_pluse(
        scalestate_0_tetw_pluse), .scalestate_0_dumpoff_ctr(
        scalestate_0_dumpoff_ctr), .top_code_0_pn_change(
        top_code_0_pn_change), .scalestate_0_dump_sustain_ctrl(
        scalestate_0_dump_sustain_ctrl), .scalestate_0_dds_conf(
        scalestate_0_dds_conf), .calcuinter_c(calcuinter_c), 
        .scalestate_0_off_test(scalestate_0_off_test), 
        .scalestate_0_load_out(scalestate_0_load_out), 
        .scalestate_0_pn_out(scalestate_0_pn_out), 
        .scalestate_0_sw_acq1(scalestate_0_sw_acq1), 
        .scalestate_0_sw_acq2(scalestate_0_sw_acq2), 
        .top_code_0_scaleload(top_code_0_scaleload), 
        .timer_top_0_clk_en_scale_0(timer_top_0_clk_en_scale_0), 
        .top_code_0_scale_rst(top_code_0_scale_rst), .GLA(GLA_net_1));
    NOR2A \xd_pad_RNIG8Q8[9]  (.A(\xd_in[9] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[9] ));
    OUTBUF ddsreset_pad (.D(ddsreset_c), .PAD(ddsreset));
    INBUF \ADC_pad[11]  (.PAD(ADC[11]), .Y(\ADC_c[11] ));
    NOR2A \xd_pad_RNITPFD[15]  (.A(\xd_in[15] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[15] ));
    NOR2A \xd_pad_RNIC8Q8[5]  (.A(\xd_in[5] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[5] ));
    topctrlchange topctrlchange_0 (.change({\change[1] , \change[0] }), 
        .GLA(GLA_net_1), .plusestate_0_sw_acq1(plusestate_0_sw_acq1), 
        .scalestate_0_sw_acq1(scalestate_0_sw_acq1), 
        .plusestate_0_state_over_n(plusestate_0_state_over_n), 
        .scalestate_0_tetw_pluse(scalestate_0_tetw_pluse), 
        .nsctrl_choice_0_intertodsp(nsctrl_choice_0_intertodsp), 
        .scalestate_0_sw_acq2(scalestate_0_sw_acq2), 
        .nsctrl_choice_0_sw_acq2(nsctrl_choice_0_sw_acq2), 
        .plusestate_0_soft_d(plusestate_0_soft_d), 
        .scalestate_0_soft_d(scalestate_0_soft_d), 
        .nsctrl_choice_0_soft_d(nsctrl_choice_0_soft_d), 
        .scalestate_0_rt_sw(scalestate_0_rt_sw), 
        .nsctrl_choice_0_rt_sw(nsctrl_choice_0_rt_sw), .net_27(net_27), 
        .rt_sw_net_1(rt_sw_net_1), .soft_dump_net_1(soft_dump_net_1), 
        .sw_acq1_c(sw_acq1_c), .sw_acq2_c(sw_acq2_c), .un1_change_2(
        \dds_change_0.un1_change_2 ), .interupt_c(interupt_c));
    BUFF \xa_pad_RNI0QR1[7]  (.A(\xa_c[7] ), .Y(\xa_c_0[7] ));
    GPMI GPMI_0 (.GPMI_VCC(VCC), .xd_1(\GPMI_0.tri_state_0.xd_1 ), 
        .tri_ctrl_c(tri_ctrl_c), .zcs2_c(zcs2_c), .net_27(net_27), 
        .xwe_c(xwe_c), .GPMI_0_code_en(GPMI_0_code_en), .GLA(GLA_net_1)
        , .gpio_c(gpio_c));
    OR3 OR3_0 (.A(DUMP_OFF_1_dump_off), .B(DUMP_OFF_0_dump_off), .C(
        DUMP_0_dump_off), .Y(dumpoff_c));
    NOR2A \xd_pad_RNI88Q8[1]  (.A(\xd_in[1] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1_0[1] ));
    plusestate plusestate_0 (.timecount_1_1({\timecount_1_1[15] , 
        \timecount_1_1[14] , \timecount_1_1[13] , \timecount_1_1[12] , 
        \timecount_1_1[11] , \timecount_1_1[10] , \timecount_1_1[9] , 
        \timecount_1_1[8] , \timecount_1_1[7] , \timecount_1_1[6] , 
        \timecount_1_1[5] , \timecount_1_1[4] , \timecount_1_1[3] , 
        \timecount_1_1[2] , \timecount_1_1[1] , \timecount_1_1[0] }), 
        .plusedata({\plusedata[15] , \plusedata[14] , \plusedata[13] , 
        \plusedata[12] , \plusedata[11] , \plusedata[10] , 
        \plusedata[9] , \plusedata[8] , \plusedata[7] , \plusedata[6] , 
        \plusedata[5] , \plusedata[4] , \plusedata[3] , \plusedata[2] , 
        \plusedata[1] , \plusedata[0] }), .GLA(GLA_net_1), 
        .plusestate_0_off_test(plusestate_0_off_test), 
        .plusestate_0_sw_acq1(plusestate_0_sw_acq1), 
        .plusestate_0_pluse_acq(plusestate_0_pluse_acq), 
        .plusestate_0_dds_config(plusestate_0_dds_config), 
        .plusestate_0_state_over_n(plusestate_0_state_over_n), 
        .top_code_0_pluse_rst(top_code_0_pluse_rst), 
        .top_code_0_pluse_lc(top_code_0_pluse_lc), 
        .top_code_0_pluseload(top_code_0_pluseload), 
        .plusestate_0_tetw_pluse(plusestate_0_tetw_pluse), 
        .timer_top_0_clk_en_pluse(timer_top_0_clk_en_pluse), 
        .plusestate_0_soft_d(plusestate_0_soft_d), 
        .top_code_0_pluse_rst_0(top_code_0_pluse_rst_0));
    bridge_div bridge_div_0 (.scaleddsdiv({\scaleddsdiv[5] , 
        \scaleddsdiv[4] , \scaleddsdiv[3] , \scaleddsdiv[2] , 
        \scaleddsdiv[1] , \scaleddsdiv[0] }), .top_code_0_bridge_load(
        top_code_0_bridge_load), .GLA(GLA_net_1), 
        .bri_dump_sw_0_reset_out(bri_dump_sw_0_reset_out), 
        .ddsclkout_c(ddsclkout_c), .clk_4f_en(clk_4f_en), 
        .pd_pulse_en_c(pd_pulse_en_c));
    OUTBUF \relayclose_on_pad[12]  (.D(\relayclose_on_c[12] ), .PAD(
        relayclose_on[12]));
    INBUF \ADC_pad[7]  (.PAD(ADC[7]), .Y(\ADC_c[7] ));
    s_acq_change s_acq_change_0 (.s_acqnum_1({\s_acqnum_1[11] , 
        \s_acqnum_1[10] , \s_acqnum_1[9] , \s_acqnum_1[8] , 
        \s_acqnum_1[7] , \s_acqnum_1[6] , \s_acqnum_1[5] , 
        \s_acqnum_1[4] , \s_acqnum_1[3] , \s_acqnum_1[2] , 
        \s_acqnum_1[1] , \s_acqnum_1[0] }), .s_acqnum_0({
        \s_acqnum_0[15] , \s_acqnum_0[14] , \s_acqnum_0[13] , 
        \s_acqnum_0[12] , \s_acqnum_0[11] , \s_acqnum_0[10] , 
        \s_acqnum_0[9] , \s_acqnum_0[8] , \s_acqnum_0[7] , 
        \s_acqnum_0[6] , \s_acqnum_0[5] , \s_acqnum_0[4] , 
        \s_acqnum_0[3] , \s_acqnum_0[2] , \s_acqnum_0[1] , 
        \s_acqnum_0[0] }), .strippluse({\strippluse[11] , 
        \strippluse[10] , \strippluse[9] , \strippluse[8] , 
        \strippluse[7] , \strippluse[6] , \strippluse[5] , 
        \strippluse[4] , \strippluse[3] , \strippluse[2] , 
        \strippluse[1] , \strippluse[0] }), .change({\change[1] , 
        \change[0] }), .s_acqnum({\s_acqnum[15] , \s_acqnum[14] , 
        \s_acqnum[13] , \s_acqnum[12] , \s_acqnum[11] , \s_acqnum[10] , 
        \s_acqnum[9] , \s_acqnum[8] , \s_acqnum[7] , \s_acqnum[6] , 
        \s_acqnum[5] , \s_acqnum[4] , \s_acqnum[3] , \s_acqnum[2] , 
        \s_acqnum[1] , \s_acqnum[0] }), .s_stripnum({\s_stripnum[11] , 
        \s_stripnum[10] , \s_stripnum[9] , \s_stripnum[8] , 
        \s_stripnum[7] , \s_stripnum[6] , \s_stripnum[5] , 
        \s_stripnum[4] , \s_stripnum[3] , \s_stripnum[2] , 
        \s_stripnum[1] , \s_stripnum[0] }), .un1_top_code_0_3_0({
        \un1_top_code_0_3_0[1] , \un1_top_code_0_3_0[0] }), 
        .s_acq_change_0_s_load(s_acq_change_0_s_load), 
        .scalestate_0_load_out(scalestate_0_load_out), 
        .top_code_0_s_load(top_code_0_s_load), .net_45(net_45), 
        .net_33_0(net_33_0), .net_27(net_27), .s_acq_change_0_s_rst(
        s_acq_change_0_s_rst), .GLA(GLA_net_1), 
        .s_acq_change_0_s_load_0(s_acq_change_0_s_load_0));
    INBUF \xa_pad[1]  (.PAD(xa[1]), .Y(\xa_c[1] ));
    BIBUF \xd_pad[14]  (.PAD(xd[14]), .D(\dataout_0[14] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[14] ));
    NOR2A \xd_pad_RNI98Q8[2]  (.A(\xd_in[2] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1_0[2] ));
    OR2 OR2_1 (.A(nsctrl_choice_0_dumpon_ctr), .B(
        dump_sustain_timer_0_start), .Y(OR2_1_Y));
    INBUF \xa_pad[3]  (.PAD(xa[3]), .Y(\xa_c[3] ));
    OUTBUF pulse_start_pad (.D(pulse_start_c), .PAD(pulse_start));
    NOR2A \xd_pad_RNIP9FD[11]  (.A(\xd_in[11] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[11] ));
    GND GND_i_0 (.Y(GND_0));
    DUMP DUMP_0 (.dumpdata({\dumpdata[11] , \dumpdata[10] , 
        \dumpdata[9] , \dumpdata[8] , \dumpdata[7] , \dumpdata[6] , 
        \dumpdata[5] , \dumpdata[4] , \dumpdata[3] , \dumpdata[2] , 
        \dumpdata[1] , \dumpdata[0] }), .dump_cho({\dump_cho[2] , 
        \dump_cho[1] , \dump_cho[0] }), .state1ms_choice_0_dump_start(
        state1ms_choice_0_dump_start), .top_code_0_dumpload(
        top_code_0_dumpload), .state1ms_choice_0_bri_cycle(
        state1ms_choice_0_bri_cycle), .bri_div_start_0(bri_div_start_0)
        , .DUMP_0_dump_off(DUMP_0_dump_off), .DUMP_0_dump_on(
        DUMP_0_dump_on), .state1ms_choice_0_reset_out(
        state1ms_choice_0_reset_out), .GLA(GLA_net_1));
    ClockManagement ClockManagement_0 (.sigtimedata({\sigtimedata[15] , 
        \sigtimedata[14] , \sigtimedata[13] , \sigtimedata[12] , 
        \sigtimedata[11] , \sigtimedata[10] , \sigtimedata[9] , 
        \sigtimedata[8] , \sigtimedata[7] , \sigtimedata[6] , 
        \sigtimedata[5] , \sigtimedata[4] , \sigtimedata[3] , 
        \sigtimedata[2] , \sigtimedata[1] , \sigtimedata[0] }), 
        .OCX40MHz_c(OCX40MHz_c), .ClockManagement_GND(GND), 
        .ClockManagement_VCC(VCC), .net_27(net_27), .clk_5K(clk_5K), 
        .sigtimeup_c(sigtimeup_c), .top_code_0_sigrst(
        top_code_0_sigrst), .GLA(GLA_net_1));
    pd_pluse_top pd_pluse_top_0 (.i_4_0(\i_4[1] ), .pd_pluse_choice({
        \pd_pluse_choice[3] , \pd_pluse_choice[2] , 
        \pd_pluse_choice[1] , \pd_pluse_choice[0] }), .i_0_0({
        \i_0_0[1] }), .pd_pluse_data({\pd_pluse_data[15] , 
        \pd_pluse_data[14] , \pd_pluse_data[13] , \pd_pluse_data[12] , 
        \pd_pluse_data[11] , \pd_pluse_data[10] , \pd_pluse_data[9] , 
        \pd_pluse_data[8] , \pd_pluse_data[7] , \pd_pluse_data[6] , 
        \pd_pluse_data[5] , \pd_pluse_data[4] , \pd_pluse_data[3] , 
        \pd_pluse_data[2] , \pd_pluse_data[1] , \pd_pluse_data[0] }), 
        .pd_pulse_en_c(pd_pulse_en_c), .net_27(net_27), 
        .top_code_0_pd_pluse_load(top_code_0_pd_pluse_load), 
        .pulse_start_c(pulse_start_c), .net_51(net_51), 
        .bri_dump_sw_0_tetw_pluse(bri_dump_sw_0_tetw_pluse), .GLA(
        GLA_net_1), .ddsclkout_c(ddsclkout_c));
    INBUF \ADC_pad[6]  (.PAD(ADC[6]), .Y(\ADC_c[6] ));
    DUMP_ON DUMP_ON_0 (.OR2_1_Y(OR2_1_Y), .OR2_2_Y(OR2_2_Y), 
        .DUMP_ON_0_dump_on(DUMP_ON_0_dump_on), .GLA(GLA_net_1));
    INBUF \xa_pad[0]  (.PAD(xa[0]), .Y(\xa_c[0] ));
    OUTBUF Q3Q6_pad (.D(Q3Q6_c), .PAD(Q3Q6));
    AND2 AND2_0 (.A(Signal_Noise_Acq_0_acq_clk), .B(
        top_code_0_acqclken), .Y(Acq_clk_c));
    OUTBUF sd_acq_en_pad (.D(sd_acq_en_c), .PAD(sd_acq_en));
    OUTBUF \relayclose_on_pad[1]  (.D(\relayclose_on_c[1] ), .PAD(
        relayclose_on[1]));
    INBUF \xa_pad[13]  (.PAD(xa[13]), .Y(\xa_c[13] ));
    OUTBUF soft_dump_pad (.D(soft_dump_c), .PAD(soft_dump));
    nsctrl_choice nsctrl_choice_0 (.nsctrl_choice_0_dumpoff_ctr(
        nsctrl_choice_0_dumpoff_ctr), .nsctrl_choice_0_dumpon_ctr(
        nsctrl_choice_0_dumpon_ctr), .nsctrl_choice_0_dumponoff_rst(
        nsctrl_choice_0_dumponoff_rst), .nsctrl_choice_0_intertodsp(
        nsctrl_choice_0_intertodsp), .nsctrl_choice_0_rt_sw(
        nsctrl_choice_0_rt_sw), .nsctrl_choice_0_soft_d(
        nsctrl_choice_0_soft_d), .GLA(GLA_net_1), 
        .nsctrl_choice_0_sw_acq2(nsctrl_choice_0_sw_acq2), 
        .noisestate_0_sw_acq2(noisestate_0_sw_acq2), 
        .scanstate_0_sw_acq2(scanstate_0_sw_acq2), 
        .top_code_0_n_s_ctrl(top_code_0_n_s_ctrl), .noisestate_0_rt_sw(
        noisestate_0_rt_sw), .scanstate_0_rt_sw(scanstate_0_rt_sw), 
        .noisestate_0_dumpon_ctr(noisestate_0_dumpon_ctr), 
        .scanstate_0_dds_conf(scanstate_0_dds_conf), 
        .top_code_0_n_s_ctrl_1(top_code_0_n_s_ctrl_1), 
        .noisestate_0_soft_d(noisestate_0_soft_d), .scanstate_0_soft_d(
        scanstate_0_soft_d), .noisestate_0_state_over_n(
        noisestate_0_state_over_n), .scanstate_0_state_over_n(
        scanstate_0_state_over_n), .top_code_0_noise_rst_0(
        top_code_0_noise_rst_0), .net_33_0(net_33_0), 
        .top_code_0_n_s_ctrl_0(top_code_0_n_s_ctrl_0), 
        .noisestate_0_dumpoff_ctr(noisestate_0_dumpoff_ctr), 
        .scanstate_0_dumpoff_ctr(scanstate_0_dumpoff_ctr), .net_27(
        net_27));
    OUTBUF pd_pulse_en_pad (.D(pd_pulse_en_c), .PAD(pd_pulse_en));
    BIBUF \xd_pad[0]  (.PAD(xd[0]), .D(\dataout_0[0] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[0] ));
    OUTBUF ddswclk_pad (.D(ddswclk_c), .PAD(ddswclk));
    NOR2A \xd_pad_RNI98Q8_0[2]  (.A(\xd_in[2] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[2] ));
    scanstate scanstate_0 (.timecount_1_0({\timecount_1_0[15] , 
        \timecount_1_0[14] , \timecount_1_0[13] , \timecount_1_0[12] , 
        \timecount_1_0[11] , \timecount_1_0[10] , \timecount_1_0[9] , 
        \timecount_1_0[8] , \timecount_1_0[7] , \timecount_1_0[6] , 
        \timecount_1_0[5] , \timecount_1_0[4] , \timecount_1_0[3] , 
        \timecount_1_0[2] , \timecount_1_0[1] , \timecount_1_0[0] }), 
        .scandata({\scandata[15] , \scandata[14] , \scandata[13] , 
        \scandata[12] , \scandata[11] , \scandata[10] , \scandata[9] , 
        \scandata[8] , \scandata[7] , \scandata[6] , \scandata[5] , 
        \scandata[4] , \scandata[3] , \scandata[2] , \scandata[1] , 
        \scandata[0] }), .GLA(GLA_net_1), .top_code_0_scanchoice(
        top_code_0_scanchoice), .top_code_0_scanload(
        top_code_0_scanload), .scanstate_0_calctrl(scanstate_0_calctrl)
        , .scanstate_0_soft_d(scanstate_0_soft_d), 
        .scanstate_0_dds_conf(scanstate_0_dds_conf), .net_33(net_33), 
        .scanstate_0_state_over_n(scanstate_0_state_over_n), 
        .scanstate_0_s_acq(scanstate_0_s_acq), 
        .scanstate_0_dumpoff_ctr(scanstate_0_dumpoff_ctr), 
        .scanstate_0_rt_sw(scanstate_0_rt_sw), .scanstate_0_sw_acq2(
        scanstate_0_sw_acq2), .net_33_0(net_33_0), 
        .timer_top_0_clk_en_scan(timer_top_0_clk_en_scan));
    NOR2A \xd_pad_RNIA8Q8[3]  (.A(\xd_in[3] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[3] ));
    INBUF \ADC_pad[4]  (.PAD(ADC[4]), .Y(\ADC_c[4] ));
    INBUF \xa_pad[9]  (.PAD(xa[9]), .Y(\xa_c[9] ));
    BUFF \xa_pad_RNIPPR1[0]  (.A(\xa_c[0] ), .Y(\xa_c_0[0] ));
    BIBUF \xd_pad[3]  (.PAD(xd[3]), .D(\dataout_0[3] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[3] ));
    OUTBUF cal_out_pad (.D(cal_out_c), .PAD(cal_out));
    INBUF \xa_pad[12]  (.PAD(xa[12]), .Y(\xa_c[12] ));
    OUTBUF \relayclose_on_pad[6]  (.D(\relayclose_on_c[6] ), .PAD(
        relayclose_on[6]));
    DUMP_OFF_DUMP_OFF_0 DUMP_OFF_0 (.bri_dump_sw_0_dumpoff_ctr(
        bri_dump_sw_0_dumpoff_ctr), .bri_dump_sw_0_reset_out_0(
        bri_dump_sw_0_reset_out_0), .DUMP_OFF_0_dump_off(
        DUMP_OFF_0_dump_off), .GLA(GLA_net_1));
    n_pluse_acq n_acq_change_0 (.n_acq_change_0_n_acq_start(
        n_acq_change_0_n_acq_start), .n_acq_change_0_n_rst_n(
        n_acq_change_0_n_rst_n), .net_27(net_27), .noisestate_0_n_acq(
        noisestate_0_n_acq), .plusestate_0_pluse_acq(
        plusestate_0_pluse_acq), .top_code_0_pluse_noise_ctrl(
        top_code_0_pluse_noise_ctrl), .top_code_0_noise_rst_0(
        top_code_0_noise_rst_0), .top_code_0_pluse_rst(
        top_code_0_pluse_rst), .GLA(GLA_net_1), 
        .n_acq_change_0_n_rst_n_0(n_acq_change_0_n_rst_n_0));
    noisestate noisestate_0 (.timecount_1({\timecount_1[15] , 
        \timecount_1[14] , \timecount_1[13] , \timecount_1[12] , 
        \timecount_1[11] , \timecount_1[10] , \timecount_1[9] , 
        \timecount_1[8] , \timecount_1[7] , \timecount_1[6] , 
        \timecount_1[5] , \timecount_1[4] , \timecount_1[3] , 
        \timecount_1[2] , \timecount_1[1] , \timecount_1[0] }), 
        .noisedata({\noisedata[15] , \noisedata[14] , \noisedata[13] , 
        \noisedata[12] , \noisedata[11] , \noisedata[10] , 
        \noisedata[9] , \noisedata[8] , \noisedata[7] , \noisedata[6] , 
        \noisedata[5] , \noisedata[4] , \noisedata[3] , \noisedata[2] , 
        \noisedata[1] , \noisedata[0] }), .GLA(GLA_net_1), 
        .noisestate_0_soft_d(noisestate_0_soft_d), 
        .noisestate_0_sw_acq2(noisestate_0_sw_acq2), 
        .noisestate_0_rt_sw(noisestate_0_rt_sw), .noisestate_0_n_acq(
        noisestate_0_n_acq), .top_code_0_nstatechoice(
        top_code_0_nstatechoice), .top_code_0_nstateload(
        top_code_0_nstateload), .noisestate_0_dumpoff_ctr(
        noisestate_0_dumpoff_ctr), .top_code_0_noise_rst(
        top_code_0_noise_rst), .noisestate_0_dumpon_ctr(
        noisestate_0_dumpon_ctr), .noisestate_0_state_over_n(
        noisestate_0_state_over_n), .top_code_0_noise_rst_0(
        top_code_0_noise_rst_0), .timer_top_0_clk_en_noise(
        timer_top_0_clk_en_noise));
    BIBUF \xd_pad[10]  (.PAD(xd[10]), .D(\dataout_0[10] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[10] ));
    INBUF \ADC_pad[2]  (.PAD(ADC[2]), .Y(\ADC_c[2] ));
    dds_change dds_change_0 (.un1_top_code_0_3_0({
        \un1_top_code_0_3_0[1] , \un1_top_code_0_3_0[0] }), .GLA(
        GLA_net_1), .top_code_0_pluse_rst(top_code_0_pluse_rst), 
        .net_45(net_45), .net_33_0(net_33_0), .plusestate_0_dds_config(
        plusestate_0_dds_config), .scalestate_0_dds_conf(
        scalestate_0_dds_conf), .scanstate_0_dds_conf(
        scanstate_0_dds_conf), .net_27(net_27), .dds_change_0_dds_conf(
        dds_change_0_dds_conf), .un1_change_2(
        \dds_change_0.un1_change_2 ), .dds_change_0_dds_rst(
        dds_change_0_dds_rst));
    OUTBUF s_acq180_pad (.D(s_acq180_c), .PAD(s_acq180));
    INBUF \xa_pad[2]  (.PAD(xa[2]), .Y(\xa_c[2] ));
    OUTBUF \relayclose_on_pad[15]  (.D(\relayclose_on_c[15] ), .PAD(
        relayclose_on[15]));
    BIBUF \xd_pad[1]  (.PAD(xd[1]), .D(\dataout_0[1] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[1] ));
    BIBUF \xd_pad[15]  (.PAD(xd[15]), .D(\dataout_0[15] ), .E(
        \GPMI_0.tri_state_0.xd_1 ), .Y(\xd_in[15] ));
    NOR2A \xd_pad_RNI88Q8_0[1]  (.A(\xd_in[1] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[1] ));
    NOR2A \xd_pad_RNIQDFD[12]  (.A(\xd_in[12] ), .B(tri_ctrl_c), .Y(
        \un1_GPMI_0_1[12] ));
    OUTBUF Q1Q8_pad (.D(Q1Q8_c), .PAD(Q1Q8));
    OUTBUF sw_acq1_pad (.D(sw_acq1_c), .PAD(sw_acq1));
    OUTBUF \relayclose_on_pad[5]  (.D(\relayclose_on_c[5] ), .PAD(
        relayclose_on[5]));
    OUTBUF \relayclose_on_pad[3]  (.D(\relayclose_on_c[3] ), .PAD(
        relayclose_on[3]));
    
endmodule
