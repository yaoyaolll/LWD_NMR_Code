//////////////////////////////////////////////////////////////////////
// Created by Actel SmartDesign Tue Dec 07 16:39:21 2010
// Testbench Template
// This is a basic testbench that instantiates your design with basic 
// clock and reset pins connected.  If your design has special
// clock/reset or testbench driver requirements then you should 
// copy this file and modify it. 
//////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

module testbench;

parameter SYSCLK_PERIOD = 100; // 10MHz

reg SYSCLK;
reg NSYSRESET;

initial
begin
    SYSCLK = 1'b0;
    NSYSRESET = 1'b0;
end

//////////////////////////////////////////////////////////////////////
// Reset Pulse
//////////////////////////////////////////////////////////////////////
initial
begin
    #(SYSCLK_PERIOD * 10 )
        NSYSRESET = 1'b1;
end


//////////////////////////////////////////////////////////////////////
// 10MHz Clock Driver
//////////////////////////////////////////////////////////////////////
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;


//////////////////////////////////////////////////////////////////////
// Instantiate Unit Under Test:  CAL
//////////////////////////////////////////////////////////////////////
CAL CAL_0 (
    // Inputs
    .clk_sys(SYSCLK),
    .rst_n(NSYSRESET),
    .cal_start({1{1'b0}}),
    .clk_dds(SYSCLK),
    .cal_load({1{1'b0}}),
    .cal_para({6{1'b0}}),

    // Outputs
    .cal( )

    // Inouts

);

endmodule

