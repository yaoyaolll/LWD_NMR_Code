//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Jan 22 17:08:03 2021
// Version: v11.9 SP6 11.9.6.7
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// top
module top(
    // Inputs
    clk100MHz,
    // Outputs
    clk1k,
    clk5MHz
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  clk100MHz;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output clk1k;
output clk5MHz;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   clk1k_net_0;
wire   clk5MHz_net_0;
wire   clk100MHz;
wire   clk5MHz_net_1;
wire   clk1k_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   VCC_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net = 1'b1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign clk5MHz_net_1 = clk5MHz_net_0;
assign clk5MHz       = clk5MHz_net_1;
assign clk1k_net_1   = clk1k_net_0;
assign clk1k         = clk1k_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------div_fre
div_fre div_fre_0(
        // Inputs
        .clk_in ( clk5MHz_net_0 ),
        // Outputs
        .clk_5k ( clk1k_net_0 ) 
        );

//--------pll_clk
pll_clk pll_clk_0(
        // Inputs
        .POWERDOWN ( VCC_net ),
        .CLKA      ( clk100MHz ),
        // Outputs
        .LOCK      (  ),
        .GLA       ( clk5MHz_net_0 ) 
        );


endmodule
