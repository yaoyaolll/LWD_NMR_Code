library verilog;
use verilog.vl_types.all;
entity n_s_change is
    port(
        un1_signal_acq_0: in     vl_logic_vector(3 downto 0);
        dataout_0_2     : out    vl_logic;
        dataout_0_3     : out    vl_logic;
        dataout_0_1     : out    vl_logic;
        dataout_0_5     : out    vl_logic;
        dataout_0_11    : out    vl_logic;
        dataout_0_7     : out    vl_logic;
        dataout_0_8     : out    vl_logic;
        dataout_0_6     : out    vl_logic;
        dataout_0_0_d0  : out    vl_logic;
        dataout_0_10    : out    vl_logic;
        dataout_0_9     : out    vl_logic;
        dataout_0_4     : out    vl_logic;
        dataout_0_0     : out    vl_logic_vector(15 downto 12);
        addresult_RNI5DQA: in     vl_logic_vector(12 downto 12);
        addresult_RNIJE5C: in     vl_logic_vector(14 downto 14);
        addresult_RNI8MQ7: in     vl_logic_vector(14 downto 14);
        addresult_RNI7DQA: in     vl_logic_vector(14 downto 14);
        addresult       : in     vl_logic_vector(15 downto 12);
        addresult_0_0   : in     vl_logic;
        addresult_0_2   : in     vl_logic;
        un1_add_reg_4_i_0: in     vl_logic;
        un1_add_reg_4_i_2: in     vl_logic;
        addresult_5_0   : in     vl_logic;
        addresult_5_2   : in     vl_logic;
        addresult_4_0   : in     vl_logic;
        addresult_4_2   : in     vl_logic;
        MX2_RD_2_inst   : in     vl_logic;
        MX2_RD_3_inst   : in     vl_logic;
        MX2_RD_1_inst   : in     vl_logic;
        MX2_RD_5_inst   : in     vl_logic;
        N_25_i_0        : in     vl_logic;
        top_code_0_n_s_ctrl: in     vl_logic;
        MX2_RD_11_inst  : in     vl_logic;
        N_20_i_0        : in     vl_logic;
        MX2_RD_7_inst   : in     vl_logic;
        N_12_i_0        : in     vl_logic;
        s_clk_div4_0_clkout: in     vl_logic;
        signal_acq_0_Signal_acq_clk: in     vl_logic;
        Signal_Noise_Acq_0_acq_clk: out    vl_logic;
        top_code_0_n_s_ctrl_1: in     vl_logic;
        MX2_RD_8_inst   : in     vl_logic;
        N_14_i_0        : in     vl_logic;
        MX2_RD_6_inst   : in     vl_logic;
        N_27_i_0        : in     vl_logic;
        MX2_RD_0_inst   : in     vl_logic;
        MX2_RD_10_inst  : in     vl_logic;
        N_18_i_0        : in     vl_logic;
        MX2_RD_9_inst   : in     vl_logic;
        N_16_i_0        : in     vl_logic;
        MX2_RD_4_inst   : in     vl_logic;
        N_22_i_0        : in     vl_logic;
        N_89            : in     vl_logic;
        N_88            : in     vl_logic;
        N_92            : in     vl_logic;
        N_86            : in     vl_logic;
        N_87            : in     vl_logic;
        N_91            : in     vl_logic;
        N_95            : in     vl_logic;
        N_97            : in     vl_logic;
        N_99            : in     vl_logic;
        N_105           : in     vl_logic;
        N_104           : in     vl_logic;
        N_108           : in     vl_logic;
        N_107           : in     vl_logic;
        N_33            : in     vl_logic;
        N_256           : in     vl_logic;
        N_111           : in     vl_logic;
        N_255           : in     vl_logic;
        N_113           : in     vl_logic;
        N_253           : in     vl_logic;
        N_115           : in     vl_logic;
        N_251           : in     vl_logic;
        top_code_0_n_s_ctrl_0: in     vl_logic;
        N_39            : in     vl_logic
    );
end n_s_change;
