library verilog;
use verilog.vl_types.all;
entity noise_addr_noise_addr_0 is
    port(
        addr_0          : out    vl_logic_vector(11 downto 0);
        n_acq_change_0_n_rst_n: in     vl_logic;
        n_acq_change_0_n_rst_n_0: in     vl_logic;
        s_clk_div4_0_clkout: in     vl_logic
    );
end noise_addr_noise_addr_0;
