library verilog;
use verilog.vl_types.all;
entity qq_coder_qq_coder_0_1 is
    port(
        i               : out    vl_logic_vector(3 downto 1);
        i_0             : out    vl_logic_vector(0 downto 0);
        qq_para2        : in     vl_logic_vector(5 downto 0);
        qq_para3        : in     vl_logic_vector(5 downto 0);
        count           : in     vl_logic_vector(4 downto 0);
        qq_para1        : in     vl_logic_vector(3 downto 0);
        GLA             : in     vl_logic;
        down            : in     vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic
    );
end qq_coder_qq_coder_0_1;
