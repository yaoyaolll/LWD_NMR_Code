library verilog;
use verilog.vl_types.all;
entity off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0 is
    port(
        count_3         : out    vl_logic_vector(4 downto 0);
        GLA             : in     vl_logic;
        bri_dump_sw_0_reset_out_0: in     vl_logic;
        off_on_state_0_state_over: in     vl_logic;
        bri_dump_sw_0_dumpoff_ctr: in     vl_logic
    );
end off_on_timer_DUMP_0_off_on_timer_0_DUMP_0_off_on_timer_0;
