library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2 is
    port(
        addresult_RNI5DQA: out    vl_logic_vector(12 downto 12);
        addresult_RNI7DQA: out    vl_logic_vector(14 downto 14);
        addresult_5_10  : out    vl_logic;
        addresult_5_8   : out    vl_logic;
        addresult_RNIDU3E: in     vl_logic_vector(4 downto 4);
        signal_data_0_iv_i_3: out    vl_logic_vector(11 downto 4);
        signal_data_iv_0_0_10: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_10_0: out    vl_logic;
        signal_data_iv_0_10_3: out    vl_logic;
        signal_data_iv_0_10_2: out    vl_logic;
        un1_ten_choice_one_0_2_0: in     vl_logic;
        un1_ten_choice_one_0_2_2: in     vl_logic;
        un1_ten_choice_one_0_2_3: in     vl_logic;
        un1_ten_choice_one_0_2_4: in     vl_logic;
        un1_ten_choice_one_0_2_5: in     vl_logic;
        un1_ten_choice_one_0_2_7: in     vl_logic;
        un1_ten_choice_one_0_2_8: in     vl_logic;
        un1_ten_choice_one_0_2_9: in     vl_logic;
        un1_ten_choice_one_0_2_10: in     vl_logic;
        un1_ten_choice_one_0_2_6: in     vl_logic;
        un1_n_s_change_0_1: in     vl_logic_vector(2 downto 0);
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_249           : in     vl_logic;
        N_252           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_215           : in     vl_logic;
        N_210           : in     vl_logic;
        N_192           : in     vl_logic;
        N_189           : in     vl_logic;
        N_179           : in     vl_logic;
        N_147           : in     vl_logic;
        N_139           : in     vl_logic;
        N_131           : in     vl_logic;
        N_123           : in     vl_logic;
        N_155           : in     vl_logic;
        N_171           : in     vl_logic;
        N_251           : in     vl_logic;
        N_241           : in     vl_logic;
        N_238           : in     vl_logic;
        N_208           : in     vl_logic;
        N_205           : in     vl_logic;
        N_224_0         : in     vl_logic;
        N_259           : in     vl_logic;
        N_221           : in     vl_logic;
        N_224           : in     vl_logic
    );
end add_reg_add_reg_2;
