//////////////////////////////////////////////////////////////////////
// Created by Actel SmartDesign Tue Jan 13 09:09:02 2015
// Testbench Template
// This is a basic testbench that instantiates your design with basic 
// clock and reset pins connected.  If your design has special
// clock/reset or testbench driver requirements then you should 
// copy this file and modify it. 
//////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

module testbench;

parameter SYSCLK_PERIOD = 100; // 10MHz

reg SYSCLK;
reg NSYSRESET;

initial
begin
    SYSCLK = 1'b0;
    NSYSRESET = 1'b0;
end

//////////////////////////////////////////////////////////////////////
// Reset Pulse
//////////////////////////////////////////////////////////////////////
initial
begin
    #(SYSCLK_PERIOD * 10 )
        NSYSRESET = 1'b1;
end


//////////////////////////////////////////////////////////////////////
// 10MHz Clock Driver
//////////////////////////////////////////////////////////////////////
always @(SYSCLK)
    #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;


//////////////////////////////////////////////////////////////////////
// Instantiate Unit Under Test:  ClockManagement
//////////////////////////////////////////////////////////////////////
ClockManagement ClockManagement_0 (
    // Inputs
    .OCX40MHz({1{1'b0}}),
    .rst_n(NSYSRESET),
    .start({1{1'b0}}),
    .timer_para({16{1'b0}}),

    // Outputs
    .GLA( ),
    .timeup( ),
    .clock_10khz( )

    // Inouts

);

endmodule

