library verilog;
use verilog.vl_types.all;
entity add_reg_add_reg_2_7 is
    port(
        addresult_RNIVJME: in     vl_logic_vector(4 downto 4);
        signal_data_0_iv_i_2: out    vl_logic_vector(11 downto 4);
        signal_data_iv_0_0_3: out    vl_logic_vector(1 downto 1);
        signal_data_iv_0_3_0: out    vl_logic;
        signal_data_iv_0_3_3: out    vl_logic;
        signal_data_iv_0_3_2: out    vl_logic;
        ADC_c           : in     vl_logic_vector(2 downto 0);
        un1_n_s_change_0_1: in     vl_logic_vector(3 downto 2);
        un1_ten_choice_one_0_4_0: in     vl_logic;
        un1_ten_choice_one_0_4_3: in     vl_logic;
        un1_ten_choice_one_0_4_1: in     vl_logic;
        un1_ten_choice_one_0_4_4: in     vl_logic;
        un1_ten_choice_one_0_4_5: in     vl_logic;
        un1_ten_choice_one_0_4_7: in     vl_logic;
        un1_ten_choice_one_0_4_8: in     vl_logic;
        un1_ten_choice_one_0_4_9: in     vl_logic;
        un1_ten_choice_one_0_4_10: in     vl_logic;
        un1_ten_choice_one_0_4_11: in     vl_logic;
        un1_ten_choice_one_0_4_6: in     vl_logic;
        un1_add_reg_4_i_2: out    vl_logic;
        un1_add_reg_4_i_0: out    vl_logic;
        s_acq_change_0_s_rst: in     vl_logic;
        signalclkctrl_0_clk_add: in     vl_logic;
        N_218           : out    vl_logic;
        N_186           : out    vl_logic;
        N_88            : out    vl_logic;
        N_104           : out    vl_logic;
        N_249           : in     vl_logic;
        N_202           : out    vl_logic;
        N_250           : in     vl_logic;
        N_249_0         : in     vl_logic;
        N_235           : out    vl_logic;
        N_212           : in     vl_logic;
        N_211           : in     vl_logic;
        N_188           : in     vl_logic;
        N_177           : in     vl_logic;
        N_145           : in     vl_logic;
        N_137           : in     vl_logic;
        N_129           : in     vl_logic;
        N_121           : in     vl_logic;
        N_153           : in     vl_logic;
        N_169           : in     vl_logic;
        N_253           : in     vl_logic;
        N_237           : in     vl_logic;
        N_204           : in     vl_logic;
        N_220           : in     vl_logic;
        N_263           : in     vl_logic;
        top_code_0_n_s_ctrl_0: in     vl_logic;
        N_217           : in     vl_logic
    );
end add_reg_add_reg_2_7;
